library verilog;
use verilog.vl_types.all;
entity altgxb_hssi_receiver is
    generic(
        channel_num     : integer := 1;
        channel_width   : integer := 20;
        deserialization_factor: integer := 10;
        run_length      : integer := 4;
        run_length_enable: string  := "OFF";
        use_8b_10b_mode : string  := "OFF";
        use_double_data_mode: string  := "OFF";
        use_rate_match_fifo: string  := "OFF";
        rate_matching_fifo_mode: string  := "NONE";
        use_channel_align: string  := "OFF";
        use_symbol_align: string  := "ON";
        use_auto_bit_slip: string  := "ON";
        synchronization_mode: string  := "NONE";
        align_pattern   : string  := "0000000101111100";
        align_pattern_length: integer := 7;
        infiniband_invalid_code: integer := 0;
        disparity_mode  : string  := "OFF";
        clk_out_mode_reference: string  := "ON";
        cruclk_period   : integer := 5000;
        cruclk_multiplier: integer := 4;
        use_cruclk_divider: string  := "OFF";
        use_parallel_feedback: string  := "OFF";
        use_post8b10b_feedback: string  := "OFF";
        send_reverse_parallel_feedback: string  := "OFF";
        use_self_test_mode: string  := "OFF";
        self_test_mode  : integer := 0;
        use_equalizer_ctrl_signal: string  := "OFF";
        enable_dc_coupling: string  := "OFF";
        equalizer_ctrl_setting: integer := 20;
        signal_threshold_select: integer := 2;
        vco_bypass      : string  := "OFF";
        force_signal_detect: string  := "OFF";
        bandwidth_type  : string  := "LOW";
        for_engineering_sample_device: string  := "ON"
    );
    port(
        datain          : in     vl_logic;
        cruclk          : in     vl_logic;
        pllclk          : in     vl_logic;
        masterclk       : in     vl_logic;
        coreclk         : in     vl_logic;
        softreset       : in     vl_logic;
        analogreset     : in     vl_logic;
        serialfdbk      : in     vl_logic;
        slpbk           : in     vl_logic;
        bitslip         : in     vl_logic;
        enacdet         : in     vl_logic;
        we              : in     vl_logic;
        re              : in     vl_logic;
        alignstatus     : in     vl_logic;
        disablefifordin : in     vl_logic;
        disablefifowrin : in     vl_logic;
        fifordin        : in     vl_logic;
        enabledeskew    : in     vl_logic;
        fiforesetrd     : in     vl_logic;
        xgmctrlin       : in     vl_logic;
        a1a2size        : in     vl_logic;
        locktorefclk    : in     vl_logic;
        locktodata      : in     vl_logic;
        parallelfdbk    : in     vl_logic_vector(9 downto 0);
        post8b10b       : in     vl_logic_vector(9 downto 0);
        equalizerctrl   : in     vl_logic_vector(2 downto 0);
        xgmdatain       : in     vl_logic_vector(7 downto 0);
        devclrn         : in     vl_logic;
        devpor          : in     vl_logic;
        syncstatusdeskew: out    vl_logic;
        adetectdeskew   : out    vl_logic;
        rdalign         : out    vl_logic;
        xgmctrldet      : out    vl_logic;
        xgmrunningdisp  : out    vl_logic;
        xgmdatavalid    : out    vl_logic;
        fifofull        : out    vl_logic;
        fifoalmostfull  : out    vl_logic;
        fifoempty       : out    vl_logic;
        fifoalmostempty : out    vl_logic;
        disablefifordout: out    vl_logic;
        disablefifowrout: out    vl_logic;
        fifordout       : out    vl_logic;
        bisterr         : out    vl_logic;
        bistdone        : out    vl_logic;
        a1a2sizeout     : out    vl_logic_vector(1 downto 0);
        signaldetect    : out    vl_logic;
        lock            : out    vl_logic;
        freqlock        : out    vl_logic;
        rlv             : out    vl_logic;
        clkout          : out    vl_logic;
        recovclkout     : out    vl_logic;
        syncstatus      : out    vl_logic_vector(1 downto 0);
        patterndetect   : out    vl_logic_vector(1 downto 0);
        ctrldetect      : out    vl_logic_vector(1 downto 0);
        errdetect       : out    vl_logic_vector(1 downto 0);
        disperr         : out    vl_logic_vector(1 downto 0);
        dataout         : out    vl_logic_vector(19 downto 0);
        xgmdataout      : out    vl_logic_vector(7 downto 0)
    );
end altgxb_hssi_receiver;
