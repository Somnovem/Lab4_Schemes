library verilog;
use verilog.vl_types.all;
entity stratixiigx_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end stratixiigx_routing_wire;
