library verilog;
use verilog.vl_types.all;
entity hardcopyiv_hssi_tx_pma is
    generic(
        lpm_type        : string  := "hardcopyiv_hssi_tx_pma";
        analog_power    : string  := "1.5V";
        channel_number  : integer := 0;
        channel_type    : string  := "auto";
        clkin_select    : integer := 0;
        clkmux_delay    : string  := "false";
        common_mode     : string  := "0.6v";
        dprio_config_mode: integer := 0;
        enable_reverse_serial_loopback: string  := "false";
        logical_channel_address: integer := 0;
        logical_protocol_hint_0: string  := "basic";
        logical_protocol_hint_1: string  := "basic";
        logical_protocol_hint_2: string  := "basic";
        logical_protocol_hint_3: string  := "basic";
        low_speed_test_select: integer := 0;
        physical_clkin0_mapping: string  := "x1";
        physical_clkin1_mapping: string  := "x4";
        physical_clkin2_mapping: string  := "xn_top";
        physical_clkin3_mapping: string  := "xn_bottom";
        physical_clkin4_mapping: string  := "hypertransport";
        preemp_pretap   : integer := 0;
        preemp_pretap_inv: string  := "false";
        preemp_tap_1    : integer := 0;
        preemp_tap_1_a  : integer := 0;
        preemp_tap_1_b  : integer := 0;
        preemp_tap_1_c  : integer := 0;
        preemp_tap_2    : integer := 0;
        preemp_tap_2_inv: string  := "false";
        protocol_hint   : string  := "basic";
        rx_detect       : integer := 0;
        serialization_factor: integer := 8;
        slew_rate       : string  := "low";
        termination     : string  := "oct 100 ohms";
        use_external_termination: string  := "false";
        use_pclk        : string  := "false";
        use_pma_direct  : string  := "false";
        use_rx_detect   : string  := "false";
        use_ser_double_data_mode: string  := "false";
        vod_selection   : integer := 0;
        vod_selection_a : integer := 0;
        vod_selection_b : integer := 0;
        vod_selection_c : integer := 0;
        vod_selection_d : integer := 0;
        \DPRIO_CHANNEL_INTERFACE_BIT\: integer := 4
    );
    port(
        datain          : in     vl_logic_vector(63 downto 0);
        datainfull      : in     vl_logic_vector(19 downto 0);
        detectrxpowerdown: in     vl_logic;
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic_vector(299 downto 0);
        extra10gin      : in     vl_logic_vector(10 downto 0);
        fastrefclk0in   : in     vl_logic_vector(1 downto 0);
        fastrefclk1in   : in     vl_logic_vector(1 downto 0);
        fastrefclk2in   : in     vl_logic_vector(1 downto 0);
        fastrefclk3in   : in     vl_logic_vector(1 downto 0);
        fastrefclk4in   : in     vl_logic_vector(1 downto 0);
        forceelecidle   : in     vl_logic;
        pclk            : in     vl_logic_vector(4 downto 0);
        powerdn         : in     vl_logic;
        refclk0in       : in     vl_logic_vector(1 downto 0);
        refclk0inpulse  : in     vl_logic;
        refclk1in       : in     vl_logic_vector(1 downto 0);
        refclk1inpulse  : in     vl_logic;
        refclk2in       : in     vl_logic_vector(1 downto 0);
        refclk2inpulse  : in     vl_logic;
        refclk3in       : in     vl_logic_vector(1 downto 0);
        refclk3inpulse  : in     vl_logic;
        refclk4in       : in     vl_logic_vector(1 downto 0);
        refclk4inpulse  : in     vl_logic;
        revserialfdbk   : in     vl_logic;
        rxdetectclk     : in     vl_logic;
        rxdetecten      : in     vl_logic;
        txpmareset      : in     vl_logic;
        clockout        : out    vl_logic;
        dataout         : out    vl_logic;
        dftout          : out    vl_logic_vector(5 downto 0);
        dprioout        : out    vl_logic_vector(299 downto 0);
        rxdetectvalidout: out    vl_logic;
        rxfoundout      : out    vl_logic;
        seriallpbkout   : out    vl_logic
    );
end hardcopyiv_hssi_tx_pma;
