library verilog;
use verilog.vl_types.all;
entity hssi_quad is
    generic(
        operation_mode  : string  := "DUPLEX";
        loopback_mode   : string  := "NONE";
        reverse_loopback_mode: string  := "NONE";
        protocol        : string  := "NONE";
        protocol_to_mode: string  := "NONE";
        tx_transmit_protocol: string  := "NONE";
        number_of_channels: integer := 4;
        channel_width   : integer := 20;
        pll_inclock_period: integer := 20000;
        data_rate       : integer := 10;
        c_use_8b_10b_mode: string  := "OFF";
        c_use_double_data_mode: string  := "OFF";
        rx_use_double_data_mode: string  := "OFF";
        c_disparity_mode: string  := "OFF";
        c_force_disparity_mode: string  := "OFF";
        cru_inclock_period: integer := 0;
        run_length      : integer := 128;
        run_length_enable: string  := "OFF";
        c_use_channel_align: string  := "OFF";
        c_use_auto_bit_slip: string  := "ON";
        c_use_rate_match_fifo: string  := "ON";
        c_use_symbol_align: string  := "ON";
        align_pattern   : string  := "";
        align_pattern_length: integer := 0;
        infiniband_invalid_code: integer := 0;
        c_clk_out_mode_reference: string  := "ON";
        c_use_fifo_mode : string  := "ON";
        intended_device_family: string  := "ALTGXB";
        deserialization_factor: integer := 8;
        pll_mult_value  : integer := 1;
        pllclk2_divisor : integer := 2;
        cruclk_mult     : integer := 0;
        cruclk_div      : string  := "";
        pllclk_mult     : integer := 1;
        pllclk0_div     : integer := 1;
        pllclk_div_adj  : integer := 1;
        use_self_test_mode: string  := "OFF";
        self_test_mode  : integer := 0;
        use_equalizer_ctrl_signal: string  := "OFF";
        equalizer_ctrl_setting: integer := 0;
        signal_threshold_select: integer := 80;
        rx_bandwidth_type: string  := "NEW_MEDIUM";
        rx_enable_dc_coupling: string  := "OFF";
        use_vod_ctrl_signal: string  := "OFF";
        vod_ctrl_setting: integer := 1000;
        use_preemphasis_ctrl_signal: string  := "OFF";
        preemphasis_ctrl_setting: integer := 0;
        use_phase_shift : string  := "ON";
        pll_bandwidth_type: string  := "LOW";
        pll_use_dc_coupling: string  := "OFF";
        rx_ppm_setting  : integer := 1000;
        device_family   : string  := "";
        use_rx_cruclk   : string  := "OFF";
        use_rx_clkout   : string  := "OFF";
        use_rx_coreclk  : string  := "OFF";
        use_tx_coreclk  : string  := "OFF";
        instantiate_transmitter_pll: string  := "OFF";
        consider_instantiate_transmitter_pll_param: string  := "OFF";
        use_generic_fifo: string  := "OFF";
        flip_rx_out     : string  := "OFF";
        flip_tx_in      : string  := "OFF";
        add_generic_fifo_we_synch_register: string  := "OFF";
        rx_dwidth_factor: integer := 2;
        for_engineering_sample_device: string  := "ON"
    );
    port(
        inclk           : in     vl_logic;
        pll_areset      : in     vl_logic;
        rx_cruclk       : in     vl_logic;
        rx_coreclk      : in     vl_logic_vector;
        rx_in           : in     vl_logic_vector;
        rx_bitslip      : in     vl_logic_vector;
        rx_enacdet      : in     vl_logic_vector;
        rx_we           : in     vl_logic_vector;
        rx_re           : in     vl_logic_vector;
        rx_slpbk        : in     vl_logic_vector;
        rx_a1a2size     : in     vl_logic_vector;
        rx_equalizerctrl: in     vl_logic_vector;
        rx_locktorefclk : in     vl_logic_vector;
        rx_locktodata   : in     vl_logic_vector;
        tx_in           : in     vl_logic_vector;
        tx_coreclk      : in     vl_logic_vector;
        tx_ctrlenable   : in     vl_logic_vector;
        tx_forcedisparity: in     vl_logic_vector;
        tx_srlpbk       : in     vl_logic_vector;
        tx_vodctrl      : in     vl_logic_vector;
        tx_preemphasisctrl: in     vl_logic_vector;
        txdigitalreset  : in     vl_logic_vector(3 downto 0);
        rxdigitalreset  : in     vl_logic_vector(3 downto 0);
        rxanalogreset   : in     vl_logic_vector(3 downto 0);
        pllenable       : in     vl_logic;
        pll_locked      : out    vl_logic;
        coreclk_out     : out    vl_logic;
        rx_out          : out    vl_logic_vector;
        rx_clkout       : out    vl_logic_vector;
        rx_locked       : out    vl_logic_vector;
        rx_freqlocked   : out    vl_logic_vector;
        rx_rlv          : out    vl_logic_vector;
        rx_syncstatus   : out    vl_logic_vector;
        rx_patterndetect: out    vl_logic_vector;
        rx_ctrldetect   : out    vl_logic_vector;
        rx_errdetect    : out    vl_logic_vector;
        rx_disperr      : out    vl_logic_vector;
        rx_signaldetect : out    vl_logic_vector;
        rx_fifoempty    : out    vl_logic_vector;
        rx_fifofull     : out    vl_logic_vector;
        rx_fifoalmostempty: out    vl_logic_vector;
        rx_fifoalmostfull: out    vl_logic_vector;
        rx_channelaligned: out    vl_logic;
        rx_bisterr      : out    vl_logic_vector;
        rx_bistdone     : out    vl_logic_vector;
        rx_a1a2sizeout  : out    vl_logic_vector;
        tx_out          : out    vl_logic_vector
    );
end hssi_quad;
