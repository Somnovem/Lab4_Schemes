library verilog;
use verilog.vl_types.all;
entity arriaii_hssi_cmu is
    generic(
        lpm_type        : string  := "arriaii_hssi_cmu";
        analog_test_bus_enable: string  := "false";
        auto_spd_deassert_ph_fifo_rst_count: integer := 0;
        auto_spd_phystatus_notify_count: integer := 0;
        bonded_quad_mode: string  := "none";
        bypass_bandgap  : string  := "false";
        central_test_bus_select: integer := 0;
        cmu_type        : string  := "regular";
        devaddr         : integer := 1;
        dprio_config_mode: integer := 0;
        in_xaui_mode    : string  := "false";
        num_con_align_chars_for_align: integer := 4;
        num_con_errors_for_align_loss: integer := 2;
        num_con_good_data_for_align_approach: integer := 3;
        offset_all_errors_align: string  := "false";
        pipe_auto_speed_nego_enable: string  := "false";
        pipe_freq_scale_mode: string  := "data width";
        pma_done_count  : integer := 0;
        portaddr        : integer := 1;
        rx0_auto_spd_self_switch_enable: string  := "false";
        rx0_channel_bonding: string  := "none";
        rx0_clk1_mux_select: string  := "recovered clock";
        rx0_clk2_mux_select: string  := "recovered clock";
        rx0_clk_pd_enable: string  := "false";
        rx0_ph_fifo_reg_mode: string  := "false";
        rx0_ph_fifo_reset_enable: string  := "false";
        rx0_ph_fifo_user_ctrl_enable: string  := "false";
        rx0_phfifo_wait_cnt: integer := 0;
        rx0_rd_clk_mux_select: string  := "int clock";
        rx0_recovered_clk_mux_select: string  := "recovered clock";
        rx0_reset_clock_output_during_digital_reset: string  := "false";
        rx0_use_double_data_mode: string  := "false";
        rx_master_direction: string  := "none";
        rx_xaui_sm_backward_compatible_enable: string  := "false";
        test_mode       : string  := "false";
        tx0_auto_spd_self_switch_enable: string  := "false";
        tx0_channel_bonding: string  := "none";
        tx0_clk_pd_enable: string  := "false";
        tx0_ph_fifo_reg_mode: string  := "false";
        tx0_ph_fifo_reset_enable: string  := "false";
        tx0_ph_fifo_user_ctrl_enable: string  := "false";
        tx0_rd_clk_mux_select: string  := "int clock";
        tx0_reset_clock_output_during_digital_reset: string  := "false";
        tx0_use_double_data_mode: string  := "false";
        tx0_wr_clk_mux_select: string  := "int_clk";
        tx_master_direction: string  := "none";
        tx_pll0_used_as_rx_cdr: string  := "false";
        tx_pll1_used_as_rx_cdr: string  := "false";
        tx_xaui_sm_backward_compatible_enable: string  := "false";
        use_deskew_fifo : string  := "false";
        vcceh_voltage   : string  := "3.0V";
        migrated_from_prev_family: string  := "false";
        protocol_hint   : string  := "basic";
        vcceh_voltage_user_specified_auto: string  := "true";
        clkdiv0_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv0_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv1_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv1_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv2_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv2_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv3_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv3_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv4_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv4_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv5_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv5_inclk1_logical_to_physical_mapping: string  := "pll1";
        cmu_divider0_inclk0_physical_mapping: string  := "pll0";
        cmu_divider0_inclk1_physical_mapping: string  := "pll1";
        cmu_divider0_inclk2_physical_mapping: string  := "x4";
        cmu_divider0_inclk3_physical_mapping: string  := "xn_t";
        cmu_divider0_inclk4_physical_mapping: string  := "xn_b";
        cmu_divider1_inclk0_physical_mapping: string  := "pll0";
        cmu_divider1_inclk1_physical_mapping: string  := "pll1";
        cmu_divider1_inclk2_physical_mapping: string  := "x4";
        cmu_divider1_inclk3_physical_mapping: string  := "xn_t";
        cmu_divider1_inclk4_physical_mapping: string  := "xn_b";
        cmu_divider2_inclk0_physical_mapping: string  := "pll0";
        cmu_divider2_inclk1_physical_mapping: string  := "pll1";
        cmu_divider2_inclk2_physical_mapping: string  := "x4";
        cmu_divider2_inclk3_physical_mapping: string  := "xn_t";
        cmu_divider2_inclk4_physical_mapping: string  := "xn_b";
        cmu_divider3_inclk0_physical_mapping: string  := "pll0";
        cmu_divider3_inclk1_physical_mapping: string  := "pll1";
        cmu_divider3_inclk2_physical_mapping: string  := "x4";
        cmu_divider3_inclk3_physical_mapping: string  := "xn_t";
        cmu_divider3_inclk4_physical_mapping: string  := "xn_b";
        cmu_divider4_inclk0_physical_mapping: string  := "pll0";
        cmu_divider4_inclk1_physical_mapping: string  := "pll1";
        cmu_divider4_inclk2_physical_mapping: string  := "x4";
        cmu_divider4_inclk3_physical_mapping: string  := "xn_t";
        cmu_divider4_inclk4_physical_mapping: string  := "xn_b";
        cmu_divider5_inclk0_physical_mapping: string  := "pll0";
        cmu_divider5_inclk1_physical_mapping: string  := "pll1";
        cmu_divider5_inclk2_physical_mapping: string  := "x4";
        cmu_divider5_inclk3_physical_mapping: string  := "xn_t";
        cmu_divider5_inclk4_physical_mapping: string  := "xn_b";
        pll0_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll0_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll0_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll0_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll0_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll0_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll0_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll0_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll0_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll0_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll1_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll1_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll1_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll1_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll1_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll1_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll1_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll1_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll1_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll1_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll2_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll2_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll2_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll2_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll2_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll2_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll2_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll2_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll2_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll2_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll3_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll3_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll3_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll3_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll3_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll3_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll3_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll3_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll3_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll3_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll4_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll4_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll4_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll4_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll4_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll4_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll4_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll4_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll4_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll4_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll5_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll5_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll5_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll5_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll5_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll5_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll5_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll5_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll5_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll5_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll0_logical_to_physical_mapping: integer := 0;
        pll1_logical_to_physical_mapping: integer := 1;
        pll2_logical_to_physical_mapping: integer := 2;
        pll3_logical_to_physical_mapping: integer := 3;
        pll4_logical_to_physical_mapping: integer := 4;
        pll5_logical_to_physical_mapping: integer := 5;
        refclk_divider0_logical_to_physical_mapping: integer := 0;
        refclk_divider1_logical_to_physical_mapping: integer := 1;
        rx0_logical_to_physical_mapping: integer := 0;
        rx1_logical_to_physical_mapping: integer := 1;
        rx2_logical_to_physical_mapping: integer := 2;
        rx3_logical_to_physical_mapping: integer := 3;
        rx4_logical_to_physical_mapping: integer := 4;
        rx5_logical_to_physical_mapping: integer := 5;
        tx0_logical_to_physical_mapping: integer := 0;
        tx1_logical_to_physical_mapping: integer := 1;
        tx2_logical_to_physical_mapping: integer := 2;
        tx3_logical_to_physical_mapping: integer := 3;
        tx4_logical_to_physical_mapping: integer := 4;
        tx5_logical_to_physical_mapping: integer := 5;
        tx0_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx0_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx0_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx0_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx0_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx1_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx1_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx1_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx1_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx1_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx2_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx2_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx2_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx2_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx2_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx3_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx3_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx3_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx3_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx3_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx4_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx4_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx4_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx4_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx4_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx5_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx5_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx5_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx5_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx5_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        sim_dump_dprio_internal_reg_at_time: integer := 0;
        sim_dump_filename: string  := "sim_dprio_dump.txt"
    );
    port(
        adet            : in     vl_logic_vector(3 downto 0);
        cmudividerdprioin: in     vl_logic_vector(599 downto 0);
        cmuplldprioin   : in     vl_logic_vector(1799 downto 0);
        dpclk           : in     vl_logic;
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic;
        dprioload       : in     vl_logic;
        extra10gin      : in     vl_logic_vector(6 downto 0);
        fixedclk        : in     vl_logic_vector(5 downto 0);
        lccmurtestbussel: in     vl_logic_vector(2 downto 0);
        pmacramtest     : in     vl_logic;
        nonuserfromcal  : in     vl_logic;
        quadreset       : in     vl_logic;
        rateswitch      : in     vl_logic;
        rateswitchdonein: in     vl_logic;
        rdalign         : in     vl_logic_vector(3 downto 0);
        rdenablesync    : in     vl_logic;
        recovclk        : in     vl_logic;
        refclkdividerdprioin: in     vl_logic_vector(1 downto 0);
        rxanalogreset   : in     vl_logic_vector(5 downto 0);
        rxclk           : in     vl_logic;
        rxcoreclk       : in     vl_logic;
        rxctrl          : in     vl_logic_vector(3 downto 0);
        rxdatain        : in     vl_logic_vector(31 downto 0);
        rxdatavalid     : in     vl_logic_vector(3 downto 0);
        rxdigitalreset  : in     vl_logic_vector(3 downto 0);
        rxpcsdprioin    : in     vl_logic_vector(1599 downto 0);
        rxphfifordenable: in     vl_logic;
        rxphfiforeset   : in     vl_logic;
        rxphfifowrdisable: in     vl_logic;
        rxpmadprioin    : in     vl_logic_vector(1799 downto 0);
        rxpowerdown     : in     vl_logic_vector(5 downto 0);
        rxrunningdisp   : in     vl_logic_vector(3 downto 0);
        scanclk         : in     vl_logic;
        scanin          : in     vl_logic_vector(22 downto 0);
        scanmode        : in     vl_logic;
        scanshift       : in     vl_logic;
        syncstatus      : in     vl_logic_vector(3 downto 0);
        testin          : in     vl_logic_vector(9999 downto 0);
        txclk           : in     vl_logic;
        txcoreclk       : in     vl_logic;
        txctrl          : in     vl_logic_vector(3 downto 0);
        txdatain        : in     vl_logic_vector(31 downto 0);
        txdigitalreset  : in     vl_logic_vector(3 downto 0);
        txpcsdprioin    : in     vl_logic_vector(599 downto 0);
        txphfiforddisable: in     vl_logic;
        txphfiforeset   : in     vl_logic;
        txphfifowrenable: in     vl_logic;
        txpllreset      : in     vl_logic_vector(1 downto 0);
        txpmadprioin    : in     vl_logic_vector(1799 downto 0);
        alignstatus     : out    vl_logic;
        autospdx4configsel: out    vl_logic;
        autospdx4rateswitchout: out    vl_logic;
        autospdx4spdchg : out    vl_logic;
        clkdivpowerdn   : out    vl_logic_vector(1 downto 0);
        cmudividerdprioout: out    vl_logic_vector(599 downto 0);
        cmuplldprioout  : out    vl_logic_vector(1799 downto 0);
        digitaltestout  : out    vl_logic_vector(9 downto 0);
        dpriodisableout : out    vl_logic;
        dpriooe         : out    vl_logic;
        dprioout        : out    vl_logic;
        enabledeskew    : out    vl_logic;
        extra10gout     : out    vl_logic;
        fiforesetrd     : out    vl_logic;
        lccmutestbus    : out    vl_logic_vector(7 downto 0);
        phfifiox4ptrsreset: out    vl_logic;
        pllpowerdn      : out    vl_logic_vector(1 downto 0);
        pllresetout     : out    vl_logic_vector(1 downto 0);
        quadresetout    : out    vl_logic;
        refclkdividerdprioout: out    vl_logic_vector(1 downto 0);
        rxadcepowerdown : out    vl_logic_vector(3 downto 0);
        rxadceresetout  : out    vl_logic_vector(3 downto 0);
        rxanalogresetout: out    vl_logic_vector(5 downto 0);
        rxcrupowerdown  : out    vl_logic_vector(5 downto 0);
        rxcruresetout   : out    vl_logic_vector(5 downto 0);
        rxctrlout       : out    vl_logic_vector(3 downto 0);
        rxdataout       : out    vl_logic_vector(31 downto 0);
        rxdigitalresetout: out    vl_logic_vector(3 downto 0);
        rxibpowerdown   : out    vl_logic_vector(5 downto 0);
        rxpcsdprioout   : out    vl_logic_vector(1599 downto 0);
        rxphfifox4byteselout: out    vl_logic;
        rxphfifox4wrclkout: out    vl_logic;
        rxphfifox4rdenableout: out    vl_logic;
        rxphfifox4wrenableout: out    vl_logic;
        rxpmadprioout   : out    vl_logic_vector(1799 downto 0);
        scanout         : out    vl_logic_vector(22 downto 0);
        testout         : out    vl_logic_vector(6999 downto 0);
        txanalogresetout: out    vl_logic_vector(5 downto 0);
        txctrlout       : out    vl_logic_vector(3 downto 0);
        txdataout       : out    vl_logic_vector(31 downto 0);
        txdetectrxpowerdown: out    vl_logic_vector(5 downto 0);
        txdigitalresetout: out    vl_logic_vector(3 downto 0);
        txdividerpowerdown: out    vl_logic_vector(5 downto 0);
        txobpowerdown   : out    vl_logic_vector(5 downto 0);
        txpcsdprioout   : out    vl_logic_vector(599 downto 0);
        txphfifox4byteselout: out    vl_logic;
        txphfifox4rdclkout: out    vl_logic;
        txphfifox4rdenableout: out    vl_logic;
        txphfifox4wrenableout: out    vl_logic;
        txpmadprioout   : out    vl_logic_vector(1799 downto 0)
    );
end arriaii_hssi_cmu;
