library verilog;
use verilog.vl_types.all;
entity \ARRIAGX_PRIM_DFFEAS\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \ARRIAGX_PRIM_DFFEAS\;
