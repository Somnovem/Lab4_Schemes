library verilog;
use verilog.vl_types.all;
entity stratixiv_hssi_tx_digi_tx_ctrl is
    port(
        soft_reset      : in     vl_logic;
        fifo_wr_clk     : in     vl_logic;
        fifo_rd_clk     : in     vl_logic;
        refclk_b_in     : in     vl_logic;
        scan_mode       : in     vl_logic;
        rindv_tx        : in     vl_logic;
        p_rlpbk         : in     vl_logic;
        selftest_en     : in     vl_logic;
        rdwidth_tx      : in     vl_logic;
        txfifo_dis      : in     vl_logic;
        rtxfifo_urst_en : in     vl_logic;
        txfifo_urst     : in     vl_logic;
        rtxfifo_lowlatency_en: in     vl_logic;
        rtxphfifopldctl_en: in     vl_logic;
        rtx_pipe_enable : in     vl_logic;
        pld_we          : in     vl_logic;
        pld_rd_dis      : in     vl_logic;
        txd             : in     vl_logic_vector(39 downto 0);
        txd_extend      : in     vl_logic_vector(3 downto 0);
        rforce_disp     : in     vl_logic;
        tx_data_sg      : in     vl_logic_vector(31 downto 0);
        tx_control_sg   : in     vl_logic_vector(3 downto 0);
        rxd_lpbk        : in     vl_logic_vector(39 downto 0);
        redund_ctl      : in     vl_logic_vector(3 downto 0);
        txd_redun       : in     vl_logic_vector(39 downto 0);
        rforce_kchar    : in     vl_logic;
        rforce_echar    : in     vl_logic;
        rtxpcsbypass_en : in     vl_logic;
        txdetectrxloopback: in     vl_logic;
        powerdown       : in     vl_logic_vector(1 downto 0);
        revloopback     : in     vl_logic;
        txswing         : in     vl_logic;
        txdeemph        : in     vl_logic;
        txmargin        : in     vl_logic_vector(2 downto 0);
        rxpolarity      : in     vl_logic;
        polinv_rx       : in     vl_logic;
        eidleinfersel   : in     vl_logic_vector(2 downto 0);
        reset_pc_ptrs   : in     vl_logic;
        reset_pc_ptrs_centrl: in     vl_logic;
        reset_pc_ptrs_quad_up: in     vl_logic;
        reset_pc_ptrs_quad_down: in     vl_logic;
        gen2ngen1       : in     vl_logic;
        gen2ngen1_bundle: in     vl_logic;
        dis_pc_byte     : in     vl_logic;
        wr_enable_centrl: in     vl_logic;
        wr_enable_quad_up: in     vl_logic;
        wr_enable_quad_down: in     vl_logic;
        rd_enable_centrl: in     vl_logic;
        rd_enable_quad_up: in     vl_logic;
        rd_enable_quad_down: in     vl_logic;
        fifo_select_in_centrl: in     vl_logic;
        fifo_select_in_quad_up: in     vl_logic;
        fifo_select_in_quad_down: in     vl_logic;
        rauto_speed_ena : in     vl_logic;
        rfreq_sel       : in     vl_logic;
        rphfifo_regmode_tx: in     vl_logic;
        rmaster_tx      : in     vl_logic;
        rmaster_up_tx   : in     vl_logic;
        txd_extend_tc   : out    vl_logic_vector(1 downto 0);
        tx_data_tc      : out    vl_logic_vector(15 downto 0);
        tx_ctl_tc       : out    vl_logic_vector(1 downto 0);
        tx_data_9_tc    : out    vl_logic_vector(1 downto 0);
        rd_enable_sync  : out    vl_logic;
        k_det           : out    vl_logic_vector(1 downto 0);
        d21_5_eq_n      : out    vl_logic_vector(1 downto 0);
        d2_2_eq_n       : out    vl_logic_vector(1 downto 0);
        wr_enable_out   : out    vl_logic;
        rd_enable_out   : out    vl_logic;
        fifo_select_out : out    vl_logic;
        ph_fifo_full    : out    vl_logic;
        ph_fifo_empty   : out    vl_logic;
        soft_reset_wclk1: out    vl_logic;
        soft_reset_rclk1: out    vl_logic;
        pipe_electric_idle: out    vl_logic;
        txdetectrxloopback_int: out    vl_logic;
        powerdown_int   : out    vl_logic_vector(1 downto 0);
        revloopback_int : out    vl_logic;
        phfifo_txswing  : out    vl_logic;
        phfifo_txdeemph : out    vl_logic;
        phfifo_txmargin : out    vl_logic_vector(2 downto 0);
        rxpolarity_int  : out    vl_logic;
        polinv_rx_int   : out    vl_logic;
        gray_eidleinfersel: out    vl_logic_vector(2 downto 0);
        wr_enable2      : out    vl_logic;
        wptr_bin        : out    vl_logic_vector(2 downto 0);
        rd_enable2      : out    vl_logic;
        rptr_bin        : out    vl_logic_vector(2 downto 0)
    );
end stratixiv_hssi_tx_digi_tx_ctrl;
