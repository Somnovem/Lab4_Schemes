library verilog;
use verilog.vl_types.all;
entity arriaii_hssi_cmu_dprio_top is
    generic(
        clkdiv0_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv0_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv1_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv1_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv2_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv2_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv3_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv3_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv4_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv4_inclk1_logical_to_physical_mapping: string  := "pll1";
        clkdiv5_inclk0_logical_to_physical_mapping: string  := "pll0";
        clkdiv5_inclk1_logical_to_physical_mapping: string  := "pll1";
        pll0_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll0_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll0_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll0_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll0_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll0_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll0_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll0_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll0_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll0_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll1_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll1_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll1_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll1_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll1_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll1_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll1_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll1_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll1_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll1_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll2_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll2_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll2_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll2_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll2_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll2_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll2_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll2_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll2_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll2_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll3_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll3_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll3_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll3_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll3_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll3_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll3_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll3_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll3_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll3_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll4_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll4_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll4_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll4_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll4_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll4_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll4_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll4_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll4_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll4_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll5_inclk0_logical_to_physical_mapping: string  := "clkrefclk0";
        pll5_inclk1_logical_to_physical_mapping: string  := "clkrefclk1";
        pll5_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll5_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll5_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll5_inclk5_logical_to_physical_mapping: string  := "iq5";
        pll5_inclk6_logical_to_physical_mapping: string  := "iq6";
        pll5_inclk7_logical_to_physical_mapping: string  := "iq7";
        pll5_inclk8_logical_to_physical_mapping: string  := "pld_clk";
        pll5_inclk9_logical_to_physical_mapping: string  := "gpll_clk";
        pll0_logical_to_physical_mapping: integer := 0;
        pll1_logical_to_physical_mapping: integer := 1;
        pll2_logical_to_physical_mapping: integer := 2;
        pll3_logical_to_physical_mapping: integer := 3;
        pll4_logical_to_physical_mapping: integer := 4;
        pll5_logical_to_physical_mapping: integer := 5;
        refclk_divider0_logical_to_physical_mapping: integer := 0;
        refclk_divider1_logical_to_physical_mapping: integer := 1;
        rx0_logical_to_physical_mapping: integer := 0;
        rx1_logical_to_physical_mapping: integer := 1;
        rx2_logical_to_physical_mapping: integer := 2;
        rx3_logical_to_physical_mapping: integer := 3;
        rx4_logical_to_physical_mapping: integer := 4;
        rx5_logical_to_physical_mapping: integer := 5;
        tx0_logical_to_physical_mapping: integer := 0;
        tx1_logical_to_physical_mapping: integer := 1;
        tx2_logical_to_physical_mapping: integer := 2;
        tx3_logical_to_physical_mapping: integer := 3;
        tx4_logical_to_physical_mapping: integer := 4;
        tx5_logical_to_physical_mapping: integer := 5;
        tx0_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx0_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx0_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx0_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx0_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx1_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx1_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx1_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx1_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx1_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx2_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx2_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx2_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx2_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx2_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx3_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx3_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx3_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx3_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx3_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx4_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx4_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx4_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx4_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx4_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        tx5_pma_inclk0_logical_to_physical_mapping: string  := "x1";
        tx5_pma_inclk1_logical_to_physical_mapping: string  := "x4";
        tx5_pma_inclk2_logical_to_physical_mapping: string  := "xn_top";
        tx5_pma_inclk3_logical_to_physical_mapping: string  := "xn_bottom";
        tx5_pma_inclk4_logical_to_physical_mapping: string  := "hypertransport";
        sim_dump_dprio_internal_reg_at_time: integer := 0;
        sim_dump_filename: string  := "sim_dprio_dump.txt"
    );
    port(
        sync_status     : in     vl_logic_vector(3 downto 0);
        align_status    : in     vl_logic;
        mdio_in         : in     vl_logic;
        mdc             : in     vl_logic;
        port_addr       : in     vl_logic_vector(4 downto 0);
        dev_addr        : in     vl_logic_vector(4 downto 0);
        mdio_dis        : in     vl_logic;
        dprioload       : in     vl_logic;
        mdio_rst        : in     vl_logic;
        cmudividerdprioin: in     vl_logic_vector(599 downto 0);
        cmuplldprioin   : in     vl_logic_vector(1799 downto 0);
        refclkdividerdprioin: in     vl_logic_vector(1 downto 0);
        rxpcsdprioin    : in     vl_logic_vector(1599 downto 0);
        rxpmadprioin    : in     vl_logic_vector(1799 downto 0);
        txpcsdprioin    : in     vl_logic_vector(599 downto 0);
        txpmadprioin    : in     vl_logic_vector(1799 downto 0);
        cmudividerdprioout: out    vl_logic_vector(599 downto 0);
        cmuplldprioout  : out    vl_logic_vector(1799 downto 0);
        refclkdividerdprioout: out    vl_logic_vector(1 downto 0);
        rxpcsdprioout   : out    vl_logic_vector(1599 downto 0);
        rxpmadprioout   : out    vl_logic_vector(1799 downto 0);
        txpcsdprioout   : out    vl_logic_vector(599 downto 0);
        txpmadprioout   : out    vl_logic_vector(1799 downto 0);
        mdio_out        : out    vl_logic;
        data_enable_n   : out    vl_logic;
        mdio_curr_st    : out    vl_logic_vector(2 downto 0)
    );
end arriaii_hssi_cmu_dprio_top;
