library verilog;
use verilog.vl_types.all;
entity cycloneiiils_and1 is
    port(
        \Y\             : out    vl_logic;
        \IN1\           : in     vl_logic
    );
end cycloneiiils_and1;
