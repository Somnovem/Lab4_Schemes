library verilog;
use verilog.vl_types.all;
entity arriaii_hssi_pma_c_adce is
    port(
        adapt_capture   : in     vl_logic;
        adapt_done      : out    vl_logic;
        atb0            : inout  vl_logic;
        atb1            : inout  vl_logic;
        atb_0           : inout  vl_logic;
        atb_1           : inout  vl_logic;
        atben           : in     vl_logic;
        atbsel          : in     vl_logic_vector(23 downto 0);
        e_clk           : out    vl_logic;
        eqa_ctrl        : out    vl_logic;
        eqa_set         : in     vl_logic_vector(2 downto 0);
        eqb_ctrl        : out    vl_logic;
        eqb_set         : in     vl_logic_vector(2 downto 0);
        eqc_ctrl        : out    vl_logic;
        eqc_set         : in     vl_logic_vector(2 downto 0);
        eqctrlout       : out    vl_logic_vector(5 downto 0);
        eqd_ctrl        : out    vl_logic;
        eqd_set         : in     vl_logic_vector(2 downto 0);
        eqin_n          : in     vl_logic;
        eqin_p          : in     vl_logic;
        eqv_ctrl        : out    vl_logic;
        eqv_set         : in     vl_logic_vector(2 downto 0);
        fine_d2aout     : out    vl_logic;
        fixed_clk       : in     vl_logic;
        hf_adapt_done   : out    vl_logic;
        hfclk_macro     : out    vl_logic;
        hfmac_cnt0_nclr : out    vl_logic;
        hfmac_cnt2_nclr : out    vl_logic;
        ib50u_c         : inout  vl_logic;
        ib50u_t         : inout  vl_logic;
        ibrgen1         : out    vl_logic;
        ibrgen2         : out    vl_logic;
        lf_adapt_done   : out    vl_logic;
        lfclk_macro     : out    vl_logic;
        lfmac_cnt0_nclr : out    vl_logic;
        lfmac_cnt2_nclr : out    vl_logic;
        lock_lf_ovd     : in     vl_logic;
        lst             : in     vl_logic_vector(4 downto 0);
        outeqn          : inout  vl_logic;
        outeqp          : inout  vl_logic;
        r_clk           : out    vl_logic;
        radce_adapt     : in     vl_logic;
        radce_digital   : in     vl_logic_vector(9 downto 0);
        radce_hflck     : in     vl_logic_vector(14 downto 0);
        radce_lflck     : in     vl_logic_vector(14 downto 0);
        radce_pdb       : in     vl_logic;
        radce_rstb      : in     vl_logic;
        radce_vod_int   : in     vl_logic_vector(2 downto 0);
        radce_vod_lsb   : in     vl_logic;
        rbit_dc         : in     vl_logic;
        rclkdiv         : in     vl_logic_vector(3 downto 0);
        rd2a_res        : in     vl_logic_vector(1 downto 0);
        rdc_freq        : in     vl_logic_vector(1 downto 0);
        rdfe_en         : in     vl_logic;
        rf_hpf          : in     vl_logic_vector(1 downto 0);
        rf_lpf          : in     vl_logic_vector(1 downto 0);
        rgenctrlout     : out    vl_logic_vector(5 downto 0);
        rhf_os          : in     vl_logic_vector(3 downto 0);
        rhyst_hf        : in     vl_logic_vector(2 downto 0);
        rhyst_lf        : in     vl_logic_vector(2 downto 0);
        rlf_os          : in     vl_logic_vector(3 downto 0);
        rrect_adj       : in     vl_logic_vector(1 downto 0);
        rrgen_bw        : in     vl_logic_vector(1 downto 0);
        rrgen_set       : in     vl_logic_vector(2 downto 0);
        rrgen_vod       : in     vl_logic_vector(2 downto 0);
        rseq_sel        : in     vl_logic_vector(1 downto 0);
        standby         : in     vl_logic;
        tmxselan        : out    vl_logic;
        tmxselbn        : out    vl_logic;
        tmxselcn        : out    vl_logic;
        tmxseldn        : out    vl_logic;
        tmxselvn        : out    vl_logic;
        updnn_hf        : out    vl_logic;
        updnn_lf        : out    vl_logic;
        vbn             : in     vl_logic;
        vccehxqyx       : inout  vl_logic;
        vccerxqyx       : inout  vl_logic;
        vctl_quiet      : inout  vl_logic;
        vssexqyx        : inout  vl_logic
    );
end arriaii_hssi_pma_c_adce;
