library verilog;
use verilog.vl_types.all;
entity hardcopyii_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end hardcopyii_routing_wire;
