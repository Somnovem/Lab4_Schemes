library verilog;
use verilog.vl_types.all;
entity arriaii_pciehip_hip_dprio_top is
    port(
        mdc             : in     vl_logic;
        dev_addr        : in     vl_logic_vector(4 downto 0);
        port_addr       : in     vl_logic_vector(4 downto 0);
        mdio_in         : in     vl_logic;
        mdio_dis        : in     vl_logic;
        mdio_rst        : in     vl_logic;
        serial_mode     : in     vl_logic;
        ser_shift_load  : in     vl_logic;
        ser_si          : in     vl_logic;
        csr_hip_in      : in     vl_logic_vector(1759 downto 0);
        hip_base_addr   : in     vl_logic_vector(7 downto 0);
        ser_so          : out    vl_logic;
        mdio_out        : out    vl_logic;
        data_enable_n   : out    vl_logic;
        curr_state      : out    vl_logic_vector(2 downto 0);
        out_hip_ctrl_1  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_2  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_3  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_4  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_5  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_6  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_7  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_8  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_9  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_10 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_11 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_12 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_13 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_14 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_15 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_16 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_17 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_18 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_19 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_20 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_21 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_22 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_23 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_24 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_25 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_26 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_27 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_28 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_29 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_30 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_31 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_32 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_33 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_34 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_35 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_36 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_37 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_38 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_39 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_40 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_41 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_42 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_43 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_44 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_45 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_46 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_47 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_48 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_49 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_50 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_51 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_52 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_53 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_54 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_55 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_56 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_57 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_58 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_59 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_60 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_61 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_62 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_63 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_64 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_65 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_66 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_67 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_68 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_69 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_70 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_71 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_72 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_73 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_74 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_75 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_76 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_77 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_78 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_79 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_80 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_81 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_82 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_83 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_84 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_85 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_86 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_87 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_88 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_89 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_90 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_91 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_92 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_93 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_94 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_95 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_96 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_97 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_98 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_99 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_100: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_101: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_102: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_103: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_104: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_105: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_106: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_107: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_108: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_109: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_110: out    vl_logic_vector(15 downto 0)
    );
end arriaii_pciehip_hip_dprio_top;
