library verilog;
use verilog.vl_types.all;
entity stratixii_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end stratixii_routing_wire;
