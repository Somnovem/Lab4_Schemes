library verilog;
use verilog.vl_types.all;
entity \TRI\ is
    port(
        \in\            : in     vl_logic;
        oe              : in     vl_logic;
        \out\           : out    vl_logic
    );
end \TRI\;
