library verilog;
use verilog.vl_types.all;
entity arriagx_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end arriagx_routing_wire;
