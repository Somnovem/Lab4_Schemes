library verilog;
use verilog.vl_types.all;
entity altgxb is
    generic(
        operation_mode  : string  := "DUPLEX";
        loopback_mode   : string  := "NONE";
        reverse_loopback_mode: string  := "NONE";
        protocol        : string  := "NONE";
        number_of_channels: integer := 20;
        number_of_quads : integer := 1;
        channel_width   : integer := 10;
        pll_inclock_period: integer := 20000;
        data_rate       : integer := 0;
        data_rate_remainder: integer := 0;
        use_8b_10b_mode : string  := "OFF";
        use_double_data_mode: string  := "OFF";
        dwidth_factor   : integer := 2;
        disparity_mode  : string  := "OFF";
        cru_inclock_period: integer := 0;
        run_length      : integer := 128;
        run_length_enable: string  := "OFF";
        use_channel_align: string  := "OFF";
        use_auto_bit_slip: string  := "ON";
        use_symbol_align: string  := "ON";
        align_pattern   : string  := "0000000101111100";
        align_pattern_length: integer := 10;
        infiniband_invalid_code: integer := 0;
        clk_out_mode_reference: string  := "ON";
        use_rate_match_fifo: string  := "ON";
        tx_termination  : integer := 0;
        use_fifo_mode   : string  := "ON";
        for_engineering_sample_device: string  := "ON";
        intended_device_family: string  := "ALTGXB";
        force_disparity_mode: string  := "OFF";
        lpm_type        : string  := "altgxb";
        use_self_test_mode: string  := "OFF";
        self_test_mode  : integer := 0;
        allow_gxb_merging: string  := "OFF";
        use_equalizer_ctrl_signal: string  := "OFF";
        equalizer_ctrl_setting: integer := 0;
        signal_threshold_select: integer := 80;
        rx_bandwidth_type: string  := "NEW_MEDIUM";
        rx_enable_dc_coupling: string  := "OFF";
        use_vod_ctrl_signal: string  := "OFF";
        vod_ctrl_setting: integer := 1000;
        use_preemphasis_ctrl_signal: string  := "OFF";
        preemphasis_ctrl_setting: integer := 0;
        use_phase_shift : string  := "ON";
        pll_bandwidth_type: string  := "LOW";
        pll_use_dc_coupling: string  := "OFF";
        rx_ppm_setting  : integer := 1000;
        device_family   : string  := "";
        use_rx_cruclk   : string  := "OFF";
        use_rx_clkout   : string  := "OFF";
        use_rx_coreclk  : string  := "OFF";
        use_tx_coreclk  : string  := "OFF";
        instantiate_transmitter_pll: string  := "OFF";
        consider_instantiate_transmitter_pll_param: string  := "OFF";
        use_generic_fifo: string  := "OFF";
        rx_force_signal_detect: string  := "OFF";
        flip_rx_out     : string  := "OFF";
        flip_tx_in      : string  := "OFF";
        add_generic_fifo_we_synch_register: string  := "OFF";
        consider_enable_tx_8b_10b_i1i2_generation: string  := "OFF";
        enable_tx_8b_10b_i1i2_generation: string  := "OFF";
        rx_data_rate    : integer := 0;
        rx_data_rate_remainder: integer := 0
    );
    port(
        inclk           : in     vl_logic_vector;
        pll_areset      : in     vl_logic_vector;
        rx_in           : in     vl_logic_vector;
        rx_coreclk      : in     vl_logic_vector;
        rx_cruclk       : in     vl_logic_vector;
        rx_aclr         : in     vl_logic_vector;
        rx_bitslip      : in     vl_logic_vector;
        rx_enacdet      : in     vl_logic_vector;
        rx_we           : in     vl_logic_vector;
        rx_re           : in     vl_logic_vector;
        rx_slpbk        : in     vl_logic_vector;
        rx_a1a2size     : in     vl_logic_vector;
        rx_equalizerctrl: in     vl_logic_vector;
        rx_locktorefclk : in     vl_logic_vector;
        rx_locktodata   : in     vl_logic_vector;
        tx_in           : in     vl_logic_vector;
        tx_coreclk      : in     vl_logic_vector;
        tx_aclr         : in     vl_logic_vector;
        tx_ctrlenable   : in     vl_logic_vector;
        tx_forcedisparity: in     vl_logic_vector;
        tx_srlpbk       : in     vl_logic_vector;
        tx_vodctrl      : in     vl_logic_vector;
        tx_preemphasisctrl: in     vl_logic_vector;
        txdigitalreset  : in     vl_logic_vector;
        rxdigitalreset  : in     vl_logic_vector;
        rxanalogreset   : in     vl_logic_vector;
        pllenable       : in     vl_logic_vector;
        pll_locked      : out    vl_logic_vector;
        coreclk_out     : out    vl_logic_vector;
        rx_out          : out    vl_logic_vector;
        rx_clkout       : out    vl_logic_vector;
        rx_locked       : out    vl_logic_vector;
        rx_freqlocked   : out    vl_logic_vector;
        rx_rlv          : out    vl_logic_vector;
        rx_syncstatus   : out    vl_logic_vector;
        rx_patterndetect: out    vl_logic_vector;
        rx_ctrldetect   : out    vl_logic_vector;
        rx_errdetect    : out    vl_logic_vector;
        rx_disperr      : out    vl_logic_vector;
        rx_signaldetect : out    vl_logic_vector;
        rx_fifoalmostempty: out    vl_logic_vector;
        rx_fifoalmostfull: out    vl_logic_vector;
        rx_channelaligned: out    vl_logic_vector;
        rx_bisterr      : out    vl_logic_vector;
        rx_bistdone     : out    vl_logic_vector;
        rx_a1a2sizeout  : out    vl_logic_vector;
        tx_out          : out    vl_logic_vector
    );
end altgxb;
