library verilog;
use verilog.vl_types.all;
entity cycloneiv_hssi_cmu is
    generic(
        lpm_type        : string  := "cycloneiv_hssi_cmu";
        coreclk_out_gated_by_quad_reset: string  := "false";
        rx0_channel_bonding: string  := "none";
        rx0_clk1_mux_select: string  := "recovered clock";
        rx0_clk2_mux_select: string  := "recovered clock";
        rx0_clk_pd_enable: string  := "false";
        rx0_ph_fifo_reg_mode: string  := "false";
        rx0_ph_fifo_reset_enable: string  := "false";
        rx0_ph_fifo_user_ctrl_enable: string  := "false";
        rx0_rd_clk_mux_select: string  := "int clock";
        rx0_recovered_clk_mux_select: string  := "recovered clock";
        rx0_reset_clock_output_during_digital_reset: string  := "false";
        rx0_use_double_data_mode: string  := "false";
        select_refclk_dig: string  := "false";
        tx0_channel_bonding: string  := "none";
        tx0_clk_pd_enable: string  := "false";
        tx0_ph_fifo_reset_enable: string  := "false";
        tx0_ph_fifo_user_ctrl_enable: string  := "false";
        tx0_rd_clk_mux_select: string  := "local";
        tx0_reset_clock_output_during_digital_reset: string  := "false";
        tx0_use_double_data_mode: string  := "false";
        tx0_wr_clk_mux_select: string  := "int_clk";
        use_coreclk_out_post_divider: string  := "false"
    );
    port(
        dpclk           : in     vl_logic;
        dpriodisable    : in     vl_logic;
        dprioin         : in     vl_logic;
        dprioload       : in     vl_logic;
        fixedclk        : in     vl_logic_vector(3 downto 0);
        nonuserfromcal  : in     vl_logic;
        pmacramtest     : in     vl_logic;
        quadreset       : in     vl_logic;
        refclkdig       : in     vl_logic;
        rxanalogreset   : in     vl_logic_vector(3 downto 0);
        rxcoreclk       : in     vl_logic;
        rxdigitalreset  : in     vl_logic_vector(3 downto 0);
        rxphfifordenable: in     vl_logic;
        rxphfiforeset   : in     vl_logic;
        rxphfifowrdisable: in     vl_logic;
        rxpowerdown     : in     vl_logic_vector(3 downto 0);
        scanclk         : in     vl_logic;
        scanmode        : in     vl_logic;
        scanshift       : in     vl_logic;
        testin          : in     vl_logic_vector(1999 downto 0);
        txclk           : in     vl_logic;
        txcoreclk       : in     vl_logic;
        txdigitalreset  : in     vl_logic_vector(3 downto 0);
        txphfiforddisable: in     vl_logic;
        txphfiforeset   : in     vl_logic;
        txphfifowrenable: in     vl_logic;
        coreclkout      : out    vl_logic;
        digitaltestout  : out    vl_logic_vector(9 downto 0);
        dpriodisableout : out    vl_logic;
        dpriooe         : out    vl_logic;
        dprioout        : out    vl_logic;
        quadresetout    : out    vl_logic;
        refclkout       : out    vl_logic;
        rxanalogresetout: out    vl_logic_vector(3 downto 0);
        rxcrupowerdown  : out    vl_logic_vector(3 downto 0);
        rxdigitalresetout: out    vl_logic_vector(3 downto 0);
        rxibpowerdown   : out    vl_logic_vector(3 downto 0);
        rxphfifox4byteselout: out    vl_logic;
        rxphfifox4rdenableout: out    vl_logic;
        rxphfifox4wrclkout: out    vl_logic;
        rxphfifox4wrenableout: out    vl_logic;
        testout         : out    vl_logic_vector(1999 downto 0);
        txanalogresetout: out    vl_logic_vector(3 downto 0);
        txdetectrxpowerdown: out    vl_logic_vector(3 downto 0);
        txdigitalresetout: out    vl_logic_vector(3 downto 0);
        txdividerpowerdown: out    vl_logic_vector(3 downto 0);
        txobpowerdown   : out    vl_logic_vector(3 downto 0);
        txphfifox4byteselout: out    vl_logic;
        txphfifox4rdclkout: out    vl_logic;
        txphfifox4rdenableout: out    vl_logic;
        txphfifox4wrenableout: out    vl_logic
    );
end cycloneiv_hssi_cmu;
