library verilog;
use verilog.vl_types.all;
entity arriagx_hssi_tx_ctrl is
    port(
        d21_5_eq_n      : out    vl_logic_vector(1 downto 0);
        d2_2_eq_n       : out    vl_logic_vector(1 downto 0);
        dwidth          : in     vl_logic;
        fifo_rd_clk     : in     vl_logic;
        fifo_select_in_ch0: in     vl_logic;
        fifo_select_in_q0_ch0: in     vl_logic;
        fifo_select_out : out    vl_logic;
        fifo_wr_clk     : in     vl_logic;
        indv            : in     vl_logic;
        k_det           : out    vl_logic_vector(1 downto 0);
        p_rlpbk         : in     vl_logic;
        ph_fifo_empty   : out    vl_logic;
        ph_fifo_full    : out    vl_logic;
        pipe_electric_idle: out    vl_logic;
        pld_rd_dis      : in     vl_logic;
        pld_we          : in     vl_logic;
        rd_enable2      : out    vl_logic;
        rd_enable_ch0   : in     vl_logic;
        rd_enable_out   : out    vl_logic;
        rd_enable_q0_ch0: in     vl_logic;
        rd_enable_sync  : out    vl_logic;
        redund_ctl      : in     vl_logic_vector(3 downto 0);
        refclk_b_in     : in     vl_logic;
        rforce_disp     : in     vl_logic;
        rforce_echar    : in     vl_logic;
        rforce_kchar    : in     vl_logic;
        rphfifo_master_sel_tx: in     vl_logic;
        rptr_bin        : out    vl_logic_vector(2 downto 0);
        rtx_pipe_enable : in     vl_logic;
        rtxfifo_lowlatency_en: in     vl_logic;
        rtxfifo_urst_en : in     vl_logic;
        rtxphfifopldctl_en: in     vl_logic;
        rxd_lpbk        : in     vl_logic_vector(39 downto 0);
        scan_mode       : in     vl_logic;
        selftest_en     : in     vl_logic;
        soft_reset      : in     vl_logic;
        soft_reset_wclk1: out    vl_logic;
        tx_control_sg   : in     vl_logic_vector(3 downto 0);
        tx_ctl_tc       : out    vl_logic_vector(1 downto 0);
        tx_data_9_tc    : out    vl_logic_vector(1 downto 0);
        tx_data_sg      : in     vl_logic_vector(31 downto 0);
        tx_data_tc      : out    vl_logic_vector(15 downto 0);
        txd             : in     vl_logic_vector(39 downto 0);
        txd_extend      : in     vl_logic_vector(3 downto 0);
        txd_extend_tc   : out    vl_logic_vector(1 downto 0);
        txd_redun       : in     vl_logic_vector(39 downto 0);
        txfifo_dis      : in     vl_logic;
        txfifo_urst     : in     vl_logic;
        wptr_bin        : out    vl_logic_vector(2 downto 0);
        wr_enable2      : out    vl_logic;
        wr_enable_ch0   : in     vl_logic;
        wr_enable_out   : out    vl_logic;
        wr_enable_q0_ch0: in     vl_logic
    );
end arriagx_hssi_tx_ctrl;
