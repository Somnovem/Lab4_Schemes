library verilog;
use verilog.vl_types.all;
entity \LPM_HINT_EVALUATION\ is
end \LPM_HINT_EVALUATION\;
