library verilog;
use verilog.vl_types.all;
entity hardcopyiii_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end hardcopyiii_routing_wire;
