library verilog;
use verilog.vl_types.all;
entity \HARDCOPYIV_PRIM_DFFE\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \HARDCOPYIV_PRIM_DFFE\;
