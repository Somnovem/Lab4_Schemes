library verilog;
use verilog.vl_types.all;
entity stratixiigx_hssi_rx_digi is
    port(
        hard_reset      : in     vl_logic;
        rxpcs_rst       : in     vl_logic;
        rxpma_rst       : in     vl_logic;
        cmpfifourst     : in     vl_logic;
        phfifourst_rx   : in     vl_logic;
        scan_mode       : in     vl_logic;
        encdt           : in     vl_logic;
        a1a2_size       : in     vl_logic;
        bitslip         : in     vl_logic;
        rdenable_rmf    : in     vl_logic;
        wrenable_rmf    : in     vl_logic;
        pld_rx_clk      : in     vl_logic;
        polinv_rx       : in     vl_logic;
        bitloc_rev_en   : in     vl_logic;
        byte_rev_en     : in     vl_logic;
        rcvd_clk_pma    : in     vl_logic;
        pudi            : in     vl_logic_vector(19 downto 0);
        sigdetni        : in     vl_logic;
        fifo_rst_rd_qd  : in     vl_logic;
        fifo_rst_rd_gp  : in     vl_logic;
        en_dskw_qd      : in     vl_logic;
        en_dskw_gp      : in     vl_logic;
        is_lane0        : in     vl_logic;
        align_status    : in     vl_logic;
        align_status_sync_0: in     vl_logic;
        align_status_sync_2: in     vl_logic;
        disable_fifo_rd_0: in     vl_logic;
        disable_fifo_rd_2: in     vl_logic;
        disable_fifo_wr_0: in     vl_logic;
        disable_fifo_wr_2: in     vl_logic;
        rx_data_rs      : in     vl_logic_vector(7 downto 0);
        rx_control_rs   : in     vl_logic;
        rcvd_clk0_pma   : in     vl_logic;
        fifo_rd_in_comp_0: in     vl_logic;
        fifo_rd_in_comp_2: in     vl_logic;
        txlp20b         : in     vl_logic_vector(19 downto 0);
        refclk_pma      : in     vl_logic;
        tx_pma_clk      : in     vl_logic;
        fref            : in     vl_logic;
        clklow          : in     vl_logic;
        bytordpld       : in     vl_logic;
        wrdisable_rx    : in     vl_logic;
        rdenable_rx     : in     vl_logic;
        pma_testbus     : in     vl_logic_vector(7 downto 0);
        encoder_testbus : in     vl_logic_vector(9 downto 0);
        tx_ctrl_testbus : in     vl_logic_vector(9 downto 0);
        rxfifo_shared_sig_in_ch0: in     vl_logic_vector(3 downto 0);
        rxfifo_shared_sig_in_q0_ch0: in     vl_logic_vector(3 downto 0);
        rx_cru_pdb      : in     vl_logic;
        rxfifo_shared_sig_out: out    vl_logic_vector(3 downto 0);
        fifo_rd_out_comp: out    vl_logic;
        rxd             : out    vl_logic_vector(63 downto 0);
        rev_loop_data   : out    vl_logic_vector(19 downto 0);
        rx_clk          : out    vl_logic;
        bisterr         : out    vl_logic;
        cg_comma        : out    vl_logic_vector(1 downto 0);
        clk_2_b         : out    vl_logic;
        rcvd_clk_pma_b  : out    vl_logic;
        sync_status     : out    vl_logic;
        disable_fifo_rd : out    vl_logic;
        disable_fifo_wr : out    vl_logic;
        align_status_sync: out    vl_logic;
        dec_data_valid  : out    vl_logic;
        dec_data        : out    vl_logic_vector(7 downto 0);
        dec_ctl         : out    vl_logic;
        running_disp    : out    vl_logic_vector(1 downto 0);
        selftest_done   : out    vl_logic;
        selftest_err    : out    vl_logic;
        err_data        : out    vl_logic_vector(15 downto 0);
        err_ctl         : out    vl_logic_vector(1 downto 0);
        prbs_done       : out    vl_logic;
        prbs_err_lt     : out    vl_logic;
        signal_detect_out: out    vl_logic;
        align_det_sync  : out    vl_logic;
        rd_align        : out    vl_logic;
        bistdone        : out    vl_logic;
        rlv             : out    vl_logic;
        rlv_lt          : out    vl_logic;
        almost_fl_rmf   : out    vl_logic;
        full_rmf        : out    vl_logic;
        almost_mt_rmf   : out    vl_logic;
        empty_rmf       : out    vl_logic;
        freq_lock       : out    vl_logic;
        full_rx         : out    vl_logic;
        empty_rx        : out    vl_logic;
        a1a2_k1k2_flag  : out    vl_logic_vector(3 downto 0);
        byteord_flag    : out    vl_logic;
        rx_pipe_clk     : out    vl_logic;
        chnl_test_bus_out: out    vl_logic_vector(9 downto 0);
        rx_pipe_soft_reset: out    vl_logic;
        rskpsetbased    : in     vl_logic;
        rtruebac2bac    : in     vl_logic;
        ralfull         : in     vl_logic_vector(3 downto 0);
        ralempty        : in     vl_logic_vector(3 downto 0);
        rcmpfifourst    : in     vl_logic;
        rphfifourstrx   : in     vl_logic;
        rcomp_size      : in     vl_logic_vector(2 downto 0);
        rcomp_pat       : in     vl_logic_vector(39 downto 0);
        rrundisp        : in     vl_logic_vector(5 downto 0);
        rib_inv_cd      : in     vl_logic_vector(1 downto 0);
        rrlv_en         : in     vl_logic;
        rsync_sm_dis    : in     vl_logic;
        rautobtalg_dis  : in     vl_logic;
        rdis_rx_disp    : in     vl_logic;
        rmatchen        : in     vl_logic;
        rgenericfifo    : in     vl_logic;
        rendec_rx       : in     vl_logic;
        rdwidth_rx      : in     vl_logic;
        rlp20ben        : in     vl_logic;
        rrxfifo_dis     : in     vl_logic;
        rpmadwidth_rx   : in     vl_logic;
        rpma_doublewidth_rx: in     vl_logic;
        renumber        : in     vl_logic_vector(2 downto 0);
        rknumber        : in     vl_logic_vector(7 downto 0);
        renpolinv_rx    : in     vl_logic;
        rgnumber        : in     vl_logic_vector(7 downto 0);
        rclkcmpsqmd     : in     vl_logic;
        rclkcmpsq1p     : in     vl_logic_vector(19 downto 0);
        rclkcmpsq1n     : in     vl_logic_vector(19 downto 0);
        rclkcmppos      : in     vl_logic;
        rosnumber       : in     vl_logic_vector(1 downto 0);
        rosbased        : in     vl_logic;
        rkchar          : in     vl_logic;
        rcascaded_8b10b_en_rx: in     vl_logic;
        resync_badcg_en : in     vl_logic_vector(1 downto 0);
        rencdt_rising   : in     vl_logic;
        rcomp_pat_porn  : in     vl_logic;
        rprbsen_rx      : in     vl_logic;
        rprbs_clr_rslt_rx: in     vl_logic;
        rbisten_rx      : in     vl_logic;
        rbist_clr_rx    : in     vl_logic;
        rwa_6g_en       : in     vl_logic;
        rbitslip_size   : in     vl_logic_vector(1 downto 0);
        rbytord_2sym_en : in     vl_logic;
        rbysync_polinv_en: in     vl_logic;
        rbitloc_rev_en  : in     vl_logic;
        rbyte_rev_en    : in     vl_logic;
        rbyteorden      : in     vl_logic_vector(1 downto 0);
        rbytordplden    : in     vl_logic;
        rphfifopldenrx  : in     vl_logic;
        rautoinsdis     : in     vl_logic;
        rppmsel         : in     vl_logic_vector(5 downto 0);
        rforce0_freqdet : in     vl_logic;
        rforce1_freqdet : in     vl_logic;
        rbytordpat      : in     vl_logic_vector(9 downto 0);
        rbytordpad      : in     vl_logic_vector(9 downto 0);
        rforce_sig_det_pcs: in     vl_logic;
        rfreerun_rx     : in     vl_logic;
        rrcvd_clk_sel   : in     vl_logic_vector(1 downto 0);
        rclk_1_sel      : in     vl_logic_vector(1 downto 0);
        rclk_2_sel      : in     vl_logic_vector(1 downto 0);
        rrx_rd_clk_sel  : in     vl_logic;
        rall_one_dect_only: in     vl_logic;
        rtest_bus_sel   : in     vl_logic_vector(2 downto 0);
        r8b10b_dec_ibm_en: in     vl_logic_vector(1 downto 0);
        rrxfifo_lowlatency_en: in     vl_logic;
        rppm_cnt_reset  : in     vl_logic;
        sel_gp_md       : in     vl_logic;
        rclkcmpinsertpad: in     vl_logic;
        rindv_rx        : in     vl_logic;
        dskwclksel      : in     vl_logic_vector(1 downto 0);
        rdskposdisp     : in     vl_logic;
        rdskchrp        : in     vl_logic_vector(9 downto 0);
        rendec_data_sel_rx: in     vl_logic;
        rphfifo_master_sel_rx: in     vl_logic;
        rprbs_sel       : in     vl_logic_vector(2 downto 0);
        rbist_sel       : in     vl_logic_vector(1 downto 0);
        rcxpat_chnl_en  : in     vl_logic_vector(1 downto 0)
    );
end stratixiigx_hssi_rx_digi;
