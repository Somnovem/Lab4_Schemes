library verilog;
use verilog.vl_types.all;
entity \LPM_DEVICE_FAMILIES\ is
end \LPM_DEVICE_FAMILIES\;
