library verilog;
use verilog.vl_types.all;
entity arriaii_and2 is
    port(
        \IN1\           : in     vl_logic;
        \IN2\           : in     vl_logic;
        \Y\             : out    vl_logic
    );
end arriaii_and2;
