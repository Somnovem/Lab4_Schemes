library verilog;
use verilog.vl_types.all;
entity hardcopyiv_pciehip_param is
    generic(
        advanced_errors : string  := "false";
        allow_rx_valid_empty: string  := "false";
        bar0_64bit_mem_space: string  := "true";
        bar0_io_space   : string  := "false";
        bar0_prefetchable: string  := "true";
        bar0_size_mask  : integer := 32;
        bar1_64bit_mem_space: string  := "false";
        bar1_io_space   : string  := "false";
        bar1_prefetchable: string  := "false";
        bar1_size_mask  : integer := 4;
        bar2_64bit_mem_space: string  := "false";
        bar2_io_space   : string  := "false";
        bar2_prefetchable: string  := "false";
        bar2_size_mask  : integer := 4;
        bar3_64bit_mem_space: string  := "false";
        bar3_io_space   : string  := "false";
        bar3_prefetchable: string  := "false";
        bar3_size_mask  : integer := 4;
        bar4_64bit_mem_space: string  := "false";
        bar4_io_space   : string  := "false";
        bar4_prefetchable: string  := "false";
        bar4_size_mask  : integer := 4;
        bar5_64bit_mem_space: string  := "false";
        bar5_io_space   : string  := "false";
        bar5_prefetchable: string  := "false";
        bar5_size_mask  : integer := 4;
        bar_io_window_size: string  := "NONE";
        bar_prefetchable: integer := 0;
        base_address    : integer := 0;
        bridge_port_ssid_support: string  := "false";
        bridge_port_vga_enable: string  := "false";
        bypass_cdc      : string  := "false";
        bypass_tl       : string  := "false";
        class_code      : integer := 16711680;
        completion_timeout: string  := "ABCD";
        core_clk_divider: integer := 1;
        core_clk_source : string  := "PLL_FIXED_CLK";
        credit_buffer_allocation_aux: string  := "BALANCED";
        deemphasis_enable: string  := "false";
        device_address  : integer := 0;
        device_id       : integer := 1;
        device_number   : integer := 0;
        diffclock_nfts_count: integer := 128;
        disable_cdc_clk_ppm: string  := "true";
        disable_async_l2_logic: string  := "false";
        disable_link_x2_support: string  := "false";
        disable_snoop_packet: integer := 0;
        dll_active_report_support: string  := "false";
        ei_delay_powerdown_count: integer := 10;
        eie_before_nfts_count: integer := 4;
        enable_adapter_half_rate_mode: string  := "false";
        enable_ch0_pclk_out: string  := "true";
        enable_completion_timeout_disable: string  := "true";
        enable_coreclk_out_half_rate: string  := "false";
        enable_ecrc_check: string  := "true";
        enable_ecrc_gen : string  := "true";
        enable_function_msi_support: string  := "true";
        enable_function_msix_support: string  := "false";
        enable_gen2_core: string  := "true";
        enable_hip_x1_loopback: string  := "false";
        enable_l1_aspm  : string  := "false";
        enable_msi_64bit_addressing: string  := "true";
        enable_msi_masking: string  := "false";
        enable_rcv0buf_a_we: string  := "true";
        enable_rcv0buf_b_re: string  := "true";
        enable_rcv0buf_output_regs: string  := "false";
        enable_rcv1buf_a_we: string  := "true";
        enable_rcv1buf_b_re: string  := "true";
        enable_rcv1buf_output_regs: string  := "false";
        enable_retrybuf_a_we: string  := "true";
        enable_retrybuf_b_re: string  := "true";
        enable_retrybuf_ecc: string  := "false";
        enable_retrybuf_output_regs: string  := "false";
        enable_retrybuf_x8_clk_stealing: integer := 0;
        enable_rx0buf_ecc: string  := "false";
        enable_rx0buf_x8_clk_stealing: integer := 0;
        enable_rx1buf_ecc: string  := "false";
        enable_rx1buf_x8_clk_stealing: integer := 0;
        enable_rx_buffer_checking: string  := "false";
        enable_rx_ei_l0s_exit_refined: string  := "false";
        enable_rx_reordering: string  := "true";
        enable_slot_register: string  := "false";
        endpoint_l0_latency: integer := 0;
        endpoint_l1_latency: integer := 0;
        expansion_base_address_register: integer := 0;
        extend_tag_field: string  := "false";
        fc_init_timer   : integer := 1024;
        flow_control_timeout_count: integer := 200;
        flow_control_update_count: integer := 30;
        gen2_diffclock_nfts_count: integer := 255;
        gen2_lane_rate_mode: string  := "false";
        gen2_sameclock_nfts_count: integer := 255;
        hot_plug_support: integer := 0;
        iei_logic       : string  := "DISABLE";
        indicator       : integer := 7;
        l01_entry_latency: integer := 31;
        l0_exit_latency_diffclock: integer := 6;
        l0_exit_latency_sameclock: integer := 6;
        l1_exit_latency_diffclock: integer := 0;
        l1_exit_latency_sameclock: integer := 0;
        lane_mask       : integer := 240;
        low_priority_vc : integer := 0;
        max_link_width  : integer := 4;
        max_payload_size: integer := 2;
        maximum_current : integer := 0;
        migrated_from_prev_family: string  := "false";
        millisecond_cycle_count: integer := 0;
        mram_bist_settings: string  := "";
        msi_function_count: integer := 2;
        msix_pba_bir    : integer := 0;
        msix_pba_offset : integer := 0;
        msix_table_bir  : integer := 0;
        msix_table_offset: integer := 0;
        msix_table_size : integer := 0;
        no_command_completed: string  := "true";
        no_soft_reset   : string  := "false";
        pcie_mode       : string  := "SHARED_MODE";
        pme_state_enable: integer := 0;
        port_link_number: integer := 1;
        port_address    : integer := 0;
        register_pipe_signals: string  := "false";
        retry_buffer_last_active_address: integer := 4095;
        retry_buffer_memory_settings: integer := 0;
        revision_id     : integer := 1;
        rx0_adap_fifo_full_value: integer := 9;
        rx1_adap_fifo_full_value: integer := 9;
        rx_cdc_full_value: integer := 12;
        rx_idl_os_count : integer := 0;
        rx_ptr0_nonposted_dpram_max: integer := 0;
        rx_ptr0_nonposted_dpram_min: integer := 0;
        rx_ptr0_posted_dpram_max: integer := 0;
        rx_ptr0_posted_dpram_min: integer := 0;
        rx_ptr1_nonposted_dpram_max: integer := 0;
        rx_ptr1_nonposted_dpram_min: integer := 0;
        rx_ptr1_posted_dpram_max: integer := 0;
        rx_ptr1_posted_dpram_min: integer := 0;
        sameclock_nfts_count: integer := 128;
        single_rx_detect: integer := 0;
        skp_os_schedule_count: integer := 0;
        slot_number     : integer := 0;
        slot_power_limit: integer := 0;
        slot_power_scale: integer := 0;
        ssid            : integer := 0;
        ssvid           : integer := 0;
        subsystem_device_id: integer := 1;
        subsystem_vendor_id: integer := 4466;
        surprise_down_error_support: string  := "false";
        tx0_adap_fifo_full_value: integer := 11;
        tx1_adap_fifo_full_value: integer := 11;
        tx_cdc_full_value: integer := 12;
        tx_cdc_stop_dummy_full_value: integer := 11;
        use_crc_forwarding: string  := "false";
        vc0_clk_enable  : string  := "true";
        vc0_rx_buffer_memory_settings: integer := 0;
        vc0_rx_flow_ctrl_compl_data: integer := 448;
        vc0_rx_flow_ctrl_compl_header: integer := 112;
        vc0_rx_flow_ctrl_nonposted_data: integer := 0;
        vc0_rx_flow_ctrl_nonposted_header: integer := 54;
        vc0_rx_flow_ctrl_posted_data: integer := 360;
        vc0_rx_flow_ctrl_posted_header: integer := 50;
        vc1_clk_enable  : string  := "false";
        vc1_rx_buffer_memory_settings: integer := 0;
        vc1_rx_flow_ctrl_compl_data: integer := 448;
        vc1_rx_flow_ctrl_compl_header: integer := 112;
        vc1_rx_flow_ctrl_nonposted_data: integer := 0;
        vc1_rx_flow_ctrl_nonposted_header: integer := 54;
        vc1_rx_flow_ctrl_posted_data: integer := 360;
        vc1_rx_flow_ctrl_posted_header: integer := 50;
        vc_arbitration  : integer := 1;
        vc_enable       : integer := 0;
        vendor_id       : integer := 4466
    );
    port(
        test_in         : in     vl_logic;
        csr_hip_in      : out    vl_logic_vector(1759 downto 0)
    );
end hardcopyiv_pciehip_param;
