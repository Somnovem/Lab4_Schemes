library verilog;
use verilog.vl_types.all;
entity \HARDCOPYII_PRIM_DFFEAS\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \HARDCOPYII_PRIM_DFFEAS\;
