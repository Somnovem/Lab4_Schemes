library verilog;
use verilog.vl_types.all;
entity hardcopyiv_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end hardcopyiv_routing_wire;
