library verilog;
use verilog.vl_types.all;
entity stratixiv_pciehip_pciexp_top_hip is
    port(
        adrd_rcv0       : out    vl_logic_vector(10 downto 0);
        adrd_rcv1       : out    vl_logic_vector(10 downto 0);
        adrd_rpl        : out    vl_logic_vector(10 downto 0);
        adwr_rcv0       : out    vl_logic_vector(10 downto 0);
        adwr_rcv1       : out    vl_logic_vector(10 downto 0);
        adwr_rpl        : out    vl_logic_vector(10 downto 0);
        clr_rxpath      : out    vl_logic;
        core_clk        : in     vl_logic;
        core_clk_vc0    : out    vl_logic;
        core_clk_vc1    : out    vl_logic;
        core_crst       : in     vl_logic;
        core_npor       : in     vl_logic;
        core_rstn       : in     vl_logic;
        core_srst       : in     vl_logic;
        cpl_err         : in     vl_logic_vector(6 downto 0);
        cpl_pending     : in     vl_logic;
        derr_rcv0       : in     vl_logic;
        derr_rcv1       : in     vl_logic;
        din_rcv0        : out    vl_logic_vector(63 downto 0);
        din_rcv1        : out    vl_logic_vector(63 downto 0);
        din_rpl         : out    vl_logic_vector(63 downto 0);
        dl_ack_phypm    : out    vl_logic_vector(1 downto 0);
        dl_ack_req_upfc : out    vl_logic;
        dl_ack_snd_upfc : out    vl_logic;
        dl_aspm_cr0     : in     vl_logic;
        dl_comclk_reg   : in     vl_logic;
        dl_ctrl_link2   : in     vl_logic_vector(12 downto 0);
        dl_current_deemp: out    vl_logic;
        dl_current_speed: out    vl_logic_vector(1 downto 0);
        dl_data_upfc    : in     vl_logic_vector(11 downto 0);
        dl_dll_req      : out    vl_logic;
        dl_err_dll      : out    vl_logic_vector(4 downto 0);
        dl_err_phy      : out    vl_logic;
        dl_hdr_upfc     : in     vl_logic_vector(7 downto 0);
        dl_inh_dllp     : in     vl_logic;
        dl_link_auto_bdw_status: out    vl_logic;
        dl_link_bdw_mng_status: out    vl_logic;
        dl_ltssm        : out    vl_logic_vector(4 downto 0);
        dl_maxpload_dcr : in     vl_logic_vector(2 downto 0);
        dl_req_phycfg   : in     vl_logic_vector(3 downto 0);
        dl_req_phypm    : in     vl_logic_vector(3 downto 0);
        dl_req_upfc     : in     vl_logic;
        dl_req_wake     : in     vl_logic;
        dl_rpbuf_emp    : out    vl_logic;
        dl_rst_enter_comp_bit: out    vl_logic;
        dl_rst_tx_margin_field: out    vl_logic;
        dl_rx_ecrcchk   : in     vl_logic;
        dl_rx_typ_pm    : out    vl_logic_vector(2 downto 0);
        dl_rx_val_fc    : out    vl_logic;
        dl_rx_val_pm    : out    vl_logic;
        dl_snd_upfc     : in     vl_logic;
        dl_tx_ack_pm    : out    vl_logic;
        dl_tx_req_pm    : in     vl_logic;
        dl_tx_typ_pm    : in     vl_logic_vector(2 downto 0);
        dl_txcfg_extsy  : in     vl_logic;
        dl_typ_upfc     : in     vl_logic_vector(1 downto 0);
        dl_up           : out    vl_logic;
        dl_vc_ctrl      : in     vl_logic_vector(7 downto 0);
        dl_vc_status    : out    vl_logic_vector(7 downto 0);
        dl_vcid_map     : in     vl_logic_vector(23 downto 0);
        dl_vcid_upfc    : in     vl_logic_vector(2 downto 0);
        dlup_exit       : out    vl_logic;
        dout_rcv0       : in     vl_logic_vector(63 downto 0);
        dout_rcv1       : in     vl_logic_vector(63 downto 0);
        dout_rpl        : in     vl_logic_vector(63 downto 0);
        eidle_infer_sel : out    vl_logic_vector(2 downto 0);
        ev_128ns        : out    vl_logic;
        ev_1us          : out    vl_logic;
        hotrst_exit     : out    vl_logic;
        int_status      : out    vl_logic_vector(3 downto 0);
        k_bar           : in     vl_logic_vector(227 downto 0);
        k_cnt           : in     vl_logic_vector(127 downto 0);
        k_conf          : in     vl_logic_vector(383 downto 0);
        k_dev           : in     vl_logic_vector(4 downto 0);
        k_gbl_hip       : in     vl_logic_vector(63 downto 0);
        k_hip           : in     vl_logic_vector(22 downto 0);
        k_port          : in     vl_logic_vector(7 downto 0);
        k_ptr0          : in     vl_logic_vector(43 downto 0);
        k_ptr1          : in     vl_logic_vector(43 downto 0);
        k_rtry          : in     vl_logic_vector(10 downto 0);
        k_vc0           : in     vl_logic_vector(55 downto 0);
        k_vc1           : in     vl_logic_vector(55 downto 0);
        k_vc2           : in     vl_logic_vector(55 downto 0);
        k_vc3           : in     vl_logic_vector(55 downto 0);
        k_vc4           : in     vl_logic_vector(55 downto 0);
        k_vc5           : in     vl_logic_vector(55 downto 0);
        k_vc6           : in     vl_logic_vector(55 downto 0);
        k_vc7           : in     vl_logic_vector(55 downto 0);
        l2_exit         : out    vl_logic;
        lane_act        : out    vl_logic_vector(3 downto 0);
        lane_reversal_enable: out    vl_logic;
        link_up         : out    vl_logic;
        lmi_ack         : out    vl_logic;
        lmi_addr        : in     vl_logic_vector(11 downto 0);
        lmi_din         : in     vl_logic_vector(31 downto 0);
        lmi_dout        : out    vl_logic_vector(31 downto 0);
        lmi_rden        : in     vl_logic;
        lmi_wren        : in     vl_logic;
        mode            : in     vl_logic_vector(1 downto 0);
        phy_clk         : in     vl_logic;
        phy_rstn        : in     vl_logic;
        phy_srst        : in     vl_logic;
        phystatus0      : in     vl_logic;
        phystatus1      : in     vl_logic;
        phystatus2      : in     vl_logic;
        phystatus3      : in     vl_logic;
        phystatus4      : in     vl_logic;
        phystatus5      : in     vl_logic;
        phystatus6      : in     vl_logic;
        phystatus7      : in     vl_logic;
        pld_clk         : in     vl_logic;
        pld_rstn        : in     vl_logic;
        pld_srst        : in     vl_logic;
        powerdown0      : out    vl_logic_vector(1 downto 0);
        powerdown1      : out    vl_logic_vector(1 downto 0);
        powerdown2      : out    vl_logic_vector(1 downto 0);
        powerdown3      : out    vl_logic_vector(1 downto 0);
        powerdown4      : out    vl_logic_vector(1 downto 0);
        powerdown5      : out    vl_logic_vector(1 downto 0);
        powerdown6      : out    vl_logic_vector(1 downto 0);
        powerdown7      : out    vl_logic_vector(1 downto 0);
        prstn           : out    vl_logic;
        rate            : out    vl_logic;
        reset_status    : out    vl_logic;
        rx_bar_dec_vc0  : out    vl_logic_vector(7 downto 0);
        rx_bar_dec_vc1  : out    vl_logic_vector(7 downto 0);
        rx_be_vc0_0     : out    vl_logic_vector(7 downto 0);
        rx_be_vc0_1     : out    vl_logic_vector(7 downto 0);
        rx_be_vc1_0     : out    vl_logic_vector(7 downto 0);
        rx_be_vc1_1     : out    vl_logic_vector(7 downto 0);
        rx_data_vc0_0   : out    vl_logic_vector(63 downto 0);
        rx_data_vc0_1   : out    vl_logic_vector(63 downto 0);
        rx_data_vc1_0   : out    vl_logic_vector(63 downto 0);
        rx_data_vc1_1   : out    vl_logic_vector(63 downto 0);
        rx_eop_vc0_0    : out    vl_logic;
        rx_eop_vc0_1    : out    vl_logic;
        rx_eop_vc1_0    : out    vl_logic;
        rx_eop_vc1_1    : out    vl_logic;
        rx_err_vc0      : out    vl_logic;
        rx_err_vc1      : out    vl_logic;
        rx_fifo_empty_vc0: out    vl_logic;
        rx_fifo_empty_vc1: out    vl_logic;
        rx_fifo_full_vc0: out    vl_logic;
        rx_fifo_full_vc1: out    vl_logic;
        rx_fifo_rdp0    : out    vl_logic_vector(3 downto 0);
        rx_fifo_rdp1    : out    vl_logic_vector(3 downto 0);
        rx_fifo_wrp0    : out    vl_logic_vector(3 downto 0);
        rx_fifo_wrp1    : out    vl_logic_vector(3 downto 0);
        rx_mask_vc0     : in     vl_logic;
        rx_mask_vc1     : in     vl_logic;
        rx_ready_vc0    : in     vl_logic;
        rx_ready_vc1    : in     vl_logic;
        rx_sop_vc0_0    : out    vl_logic;
        rx_sop_vc0_1    : out    vl_logic;
        rx_sop_vc1_0    : out    vl_logic;
        rx_sop_vc1_1    : out    vl_logic;
        rx_valid_vc0    : out    vl_logic;
        rx_valid_vc1    : out    vl_logic;
        rxdata0         : in     vl_logic_vector(7 downto 0);
        rxdata1         : in     vl_logic_vector(7 downto 0);
        rxdata2         : in     vl_logic_vector(7 downto 0);
        rxdata3         : in     vl_logic_vector(7 downto 0);
        rxdata4         : in     vl_logic_vector(7 downto 0);
        rxdata5         : in     vl_logic_vector(7 downto 0);
        rxdata6         : in     vl_logic_vector(7 downto 0);
        rxdata7         : in     vl_logic_vector(7 downto 0);
        rxdatak0        : in     vl_logic;
        rxdatak1        : in     vl_logic;
        rxdatak2        : in     vl_logic;
        rxdatak3        : in     vl_logic;
        rxdatak4        : in     vl_logic;
        rxdatak5        : in     vl_logic;
        rxdatak6        : in     vl_logic;
        rxdatak7        : in     vl_logic;
        rxelecidle0     : in     vl_logic;
        rxelecidle1     : in     vl_logic;
        rxelecidle2     : in     vl_logic;
        rxelecidle3     : in     vl_logic;
        rxelecidle4     : in     vl_logic;
        rxelecidle5     : in     vl_logic;
        rxelecidle6     : in     vl_logic;
        rxelecidle7     : in     vl_logic;
        rxpolarity0     : out    vl_logic;
        rxpolarity1     : out    vl_logic;
        rxpolarity2     : out    vl_logic;
        rxpolarity3     : out    vl_logic;
        rxpolarity4     : out    vl_logic;
        rxpolarity5     : out    vl_logic;
        rxpolarity6     : out    vl_logic;
        rxpolarity7     : out    vl_logic;
        rxstatus0       : in     vl_logic_vector(2 downto 0);
        rxstatus1       : in     vl_logic_vector(2 downto 0);
        rxstatus2       : in     vl_logic_vector(2 downto 0);
        rxstatus3       : in     vl_logic_vector(2 downto 0);
        rxstatus4       : in     vl_logic_vector(2 downto 0);
        rxstatus5       : in     vl_logic_vector(2 downto 0);
        rxstatus6       : in     vl_logic_vector(2 downto 0);
        rxstatus7       : in     vl_logic_vector(2 downto 0);
        rxvalid0        : in     vl_logic;
        rxvalid1        : in     vl_logic;
        rxvalid2        : in     vl_logic;
        rxvalid3        : in     vl_logic;
        rxvalid4        : in     vl_logic;
        rxvalid5        : in     vl_logic;
        rxvalid6        : in     vl_logic;
        rxvalid7        : in     vl_logic;
        scan_mode       : in     vl_logic;
        serr_out        : out    vl_logic;
        successful_speed_negotiation_int: out    vl_logic;
        swdn_in         : in     vl_logic_vector(2 downto 0);
        swdn_wake       : out    vl_logic;
        swup_hotrst     : out    vl_logic;
        swup_in         : in     vl_logic_vector(6 downto 0);
        test_in_hip     : in     vl_logic_vector(31 downto 0);
        test_out_hip    : out    vl_logic_vector(63 downto 0);
        tl_aer_msi_num  : in     vl_logic_vector(4 downto 0);
        tl_app_inta_ack : out    vl_logic;
        tl_app_inta_sts : in     vl_logic;
        tl_app_msi_ack  : out    vl_logic;
        tl_app_msi_num  : in     vl_logic_vector(4 downto 0);
        tl_app_msi_req  : in     vl_logic;
        tl_app_msi_tc   : in     vl_logic_vector(2 downto 0);
        tl_cfg_add      : out    vl_logic_vector(3 downto 0);
        tl_cfg_ctl      : out    vl_logic_vector(31 downto 0);
        tl_cfg_ctl_wr   : out    vl_logic;
        tl_cfg_sts      : out    vl_logic_vector(52 downto 0);
        tl_cfg_sts_wr   : out    vl_logic;
        tl_hpg_ctrler   : in     vl_logic_vector(4 downto 0);
        tl_pex_msi_num  : in     vl_logic_vector(4 downto 0);
        tl_pm_auxpwr    : in     vl_logic;
        tl_pm_data      : in     vl_logic_vector(9 downto 0);
        tl_pm_event     : in     vl_logic;
        tl_pme_to_cr    : in     vl_logic;
        tl_pme_to_sr    : out    vl_logic;
        tl_slotclk_cfg  : in     vl_logic;
        tx_cred_vc0     : out    vl_logic_vector(35 downto 0);
        tx_cred_vc1     : out    vl_logic_vector(35 downto 0);
        tx_data_vc0_0   : in     vl_logic_vector(63 downto 0);
        tx_data_vc0_1   : in     vl_logic_vector(63 downto 0);
        tx_data_vc1_0   : in     vl_logic_vector(63 downto 0);
        tx_data_vc1_1   : in     vl_logic_vector(63 downto 0);
        tx_deemph       : out    vl_logic;
        tx_eop_vc0_0    : in     vl_logic;
        tx_eop_vc0_1    : in     vl_logic;
        tx_eop_vc1_0    : in     vl_logic;
        tx_eop_vc1_1    : in     vl_logic;
        tx_err_vc0      : in     vl_logic;
        tx_err_vc1      : in     vl_logic;
        tx_fifo_empty_vc0: out    vl_logic;
        tx_fifo_empty_vc1: out    vl_logic;
        tx_fifo_full_vc0: out    vl_logic;
        tx_fifo_full_vc1: out    vl_logic;
        tx_fifo_rdp_vc0 : out    vl_logic_vector(3 downto 0);
        tx_fifo_rdp_vc1 : out    vl_logic_vector(3 downto 0);
        tx_fifo_wrp_vc0 : out    vl_logic_vector(3 downto 0);
        tx_fifo_wrp_vc1 : out    vl_logic_vector(3 downto 0);
        tx_margin       : out    vl_logic_vector(2 downto 0);
        tx_ready_vc0    : out    vl_logic;
        tx_ready_vc1    : out    vl_logic;
        tx_sop_vc0_0    : in     vl_logic;
        tx_sop_vc0_1    : in     vl_logic;
        tx_sop_vc1_0    : in     vl_logic;
        tx_sop_vc1_1    : in     vl_logic;
        tx_valid_vc0    : in     vl_logic;
        tx_valid_vc1    : in     vl_logic;
        txcompl0        : out    vl_logic;
        txcompl1        : out    vl_logic;
        txcompl2        : out    vl_logic;
        txcompl3        : out    vl_logic;
        txcompl4        : out    vl_logic;
        txcompl5        : out    vl_logic;
        txcompl6        : out    vl_logic;
        txcompl7        : out    vl_logic;
        txdata0         : out    vl_logic_vector(7 downto 0);
        txdata1         : out    vl_logic_vector(7 downto 0);
        txdata2         : out    vl_logic_vector(7 downto 0);
        txdata3         : out    vl_logic_vector(7 downto 0);
        txdata4         : out    vl_logic_vector(7 downto 0);
        txdata5         : out    vl_logic_vector(7 downto 0);
        txdata6         : out    vl_logic_vector(7 downto 0);
        txdata7         : out    vl_logic_vector(7 downto 0);
        txdatak0        : out    vl_logic;
        txdatak1        : out    vl_logic;
        txdatak2        : out    vl_logic;
        txdatak3        : out    vl_logic;
        txdatak4        : out    vl_logic;
        txdatak5        : out    vl_logic;
        txdatak6        : out    vl_logic;
        txdatak7        : out    vl_logic;
        txdetectrx0     : out    vl_logic;
        txdetectrx1     : out    vl_logic;
        txdetectrx2     : out    vl_logic;
        txdetectrx3     : out    vl_logic;
        txdetectrx4     : out    vl_logic;
        txdetectrx5     : out    vl_logic;
        txdetectrx6     : out    vl_logic;
        txdetectrx7     : out    vl_logic;
        txelecidle0     : out    vl_logic;
        txelecidle1     : out    vl_logic;
        txelecidle2     : out    vl_logic;
        txelecidle3     : out    vl_logic;
        txelecidle4     : out    vl_logic;
        txelecidle5     : out    vl_logic;
        txelecidle6     : out    vl_logic;
        txelecidle7     : out    vl_logic;
        urstn           : out    vl_logic;
        usrst           : out    vl_logic;
        wake_oen        : out    vl_logic;
        wren_rcv0       : out    vl_logic;
        wren_rcv1       : out    vl_logic;
        wren_rpl        : out    vl_logic
    );
end stratixiv_pciehip_pciexp_top_hip;
