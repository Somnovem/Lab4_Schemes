library verilog;
use verilog.vl_types.all;
entity \ALTERA_MF_HINT_EVALUATION\ is
end \ALTERA_MF_HINT_EVALUATION\;
