library verilog;
use verilog.vl_types.all;
entity arriaii_pciehip_dprio_reg is
    port(
        mdio_rst        : in     vl_logic;
        mdio_wr         : in     vl_logic;
        reg_addr        : in     vl_logic_vector(15 downto 0);
        mdc             : in     vl_logic;
        mbus_in         : in     vl_logic_vector(15 downto 0);
        serial_mode     : in     vl_logic;
        mdio_dis        : in     vl_logic;
        ser_shift_load  : in     vl_logic;
        si              : in     vl_logic;
        ext_hip_ctrl_1  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_2  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_3  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_4  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_5  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_6  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_7  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_8  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_9  : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_10 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_11 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_12 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_13 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_14 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_15 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_16 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_17 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_18 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_19 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_20 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_21 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_22 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_23 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_24 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_25 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_26 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_27 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_28 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_29 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_30 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_31 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_32 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_33 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_34 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_35 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_36 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_37 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_38 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_39 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_40 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_41 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_42 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_43 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_44 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_45 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_46 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_47 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_48 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_49 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_50 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_51 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_52 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_53 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_54 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_55 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_56 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_57 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_58 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_59 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_60 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_61 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_62 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_63 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_64 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_65 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_66 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_67 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_68 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_69 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_70 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_71 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_72 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_73 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_74 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_75 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_76 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_77 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_78 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_79 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_80 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_81 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_82 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_83 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_84 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_85 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_86 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_87 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_88 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_89 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_90 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_91 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_92 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_93 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_94 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_95 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_96 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_97 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_98 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_99 : in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_100: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_101: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_102: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_103: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_104: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_105: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_106: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_107: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_108: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_109: in     vl_logic_vector(15 downto 0);
        ext_hip_ctrl_110: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_1: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_2: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_3: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_4: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_5: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_6: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_7: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_8: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_9: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_10: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_11: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_12: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_13: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_14: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_15: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_16: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_17: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_18: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_19: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_20: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_21: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_22: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_23: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_24: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_25: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_26: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_27: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_28: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_29: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_30: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_31: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_32: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_33: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_34: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_35: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_36: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_37: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_38: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_39: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_40: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_41: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_42: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_43: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_44: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_45: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_46: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_47: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_48: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_49: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_50: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_51: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_52: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_53: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_54: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_55: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_56: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_57: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_58: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_59: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_60: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_61: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_62: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_63: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_64: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_65: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_66: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_67: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_68: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_69: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_70: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_71: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_72: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_73: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_74: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_75: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_76: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_77: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_78: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_79: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_80: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_81: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_82: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_83: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_84: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_85: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_86: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_87: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_88: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_89: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_90: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_91: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_92: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_93: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_94: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_95: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_96: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_97: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_98: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_99: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_100: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_101: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_102: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_103: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_104: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_105: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_106: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_107: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_108: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_109: in     vl_logic_vector(15 downto 0);
        targ_addr_ctrl_110: in     vl_logic_vector(15 downto 0);
        out_hip_ctrl_1  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_2  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_3  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_4  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_5  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_6  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_7  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_8  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_9  : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_10 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_11 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_12 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_13 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_14 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_15 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_16 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_17 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_18 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_19 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_20 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_21 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_22 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_23 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_24 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_25 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_26 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_27 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_28 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_29 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_30 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_31 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_32 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_33 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_34 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_35 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_36 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_37 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_38 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_39 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_40 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_41 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_42 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_43 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_44 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_45 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_46 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_47 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_48 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_49 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_50 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_51 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_52 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_53 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_54 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_55 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_56 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_57 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_58 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_59 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_60 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_61 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_62 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_63 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_64 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_65 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_66 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_67 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_68 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_69 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_70 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_71 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_72 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_73 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_74 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_75 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_76 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_77 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_78 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_79 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_80 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_81 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_82 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_83 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_84 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_85 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_86 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_87 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_88 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_89 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_90 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_91 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_92 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_93 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_94 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_95 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_96 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_97 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_98 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_99 : out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_100: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_101: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_102: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_103: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_104: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_105: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_106: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_107: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_108: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_109: out    vl_logic_vector(15 downto 0);
        out_hip_ctrl_110: out    vl_logic_vector(15 downto 0);
        so              : out    vl_logic
    );
end arriaii_pciehip_dprio_reg;
