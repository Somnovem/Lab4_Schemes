library verilog;
use verilog.vl_types.all;
entity stratixiigx_hssi_cmu_dprio_top is
    generic(
        rx_dprio_width  : integer := 800;
        tx_dprio_width  : integer := 400;
        rx0_phy         : integer := 0;
        rx1_phy         : integer := 1;
        rx2_phy         : integer := 2;
        rx3_phy         : integer := 3;
        tx0_phy         : integer := 0;
        tx1_phy         : integer := 1;
        tx2_phy         : integer := 2;
        tx3_phy         : integer := 3;
        rx0_cru_clock0_physical_mapping: string  := "refclk0";
        rx0_cru_clock1_physical_mapping: string  := "refclk1";
        rx0_cru_clock2_physical_mapping: string  := "iq0";
        rx0_cru_clock3_physical_mapping: string  := "iq1";
        rx0_cru_clock4_physical_mapping: string  := "iq2";
        rx0_cru_clock5_physical_mapping: string  := "iq3";
        rx0_cru_clock6_physical_mapping: string  := "iq4";
        rx0_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx0_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        rx1_cru_clock0_physical_mapping: string  := "refclk0";
        rx1_cru_clock1_physical_mapping: string  := "refclk1";
        rx1_cru_clock2_physical_mapping: string  := "iq0";
        rx1_cru_clock3_physical_mapping: string  := "iq1";
        rx1_cru_clock4_physical_mapping: string  := "iq2";
        rx1_cru_clock5_physical_mapping: string  := "iq3";
        rx1_cru_clock6_physical_mapping: string  := "iq4";
        rx1_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx1_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        rx2_cru_clock0_physical_mapping: string  := "refclk0";
        rx2_cru_clock1_physical_mapping: string  := "refclk1";
        rx2_cru_clock2_physical_mapping: string  := "iq0";
        rx2_cru_clock3_physical_mapping: string  := "iq1";
        rx2_cru_clock4_physical_mapping: string  := "iq2";
        rx2_cru_clock5_physical_mapping: string  := "iq3";
        rx2_cru_clock6_physical_mapping: string  := "iq4";
        rx2_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx2_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        rx3_cru_clock0_physical_mapping: string  := "refclk0";
        rx3_cru_clock1_physical_mapping: string  := "refclk1";
        rx3_cru_clock2_physical_mapping: string  := "iq0";
        rx3_cru_clock3_physical_mapping: string  := "iq1";
        rx3_cru_clock4_physical_mapping: string  := "iq2";
        rx3_cru_clock5_physical_mapping: string  := "iq3";
        rx3_cru_clock6_physical_mapping: string  := "iq4";
        rx3_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx3_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        tx0_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx0_pll_fast_clk1_physical_mapping: string  := "pll1";
        tx1_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx1_pll_fast_clk1_physical_mapping: string  := "pll1";
        tx2_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx2_pll_fast_clk1_physical_mapping: string  := "pll1";
        tx3_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx3_pll_fast_clk1_physical_mapping: string  := "pll1";
        pll0_phy        : integer := 0;
        pll1_phy        : integer := 1;
        pll2_phy        : integer := 2;
        pll0_inclk0_logical_to_physical_mapping: string  := "iq0";
        pll0_inclk1_logical_to_physical_mapping: string  := "iq1";
        pll0_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll0_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll0_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll0_inclk5_logical_to_physical_mapping: string  := "pld_clk";
        pll0_inclk6_logical_to_physical_mapping: string  := "clkrefclk0";
        pll0_inclk7_logical_to_physical_mapping: string  := "clkrefclk1";
        pll1_inclk0_logical_to_physical_mapping: string  := "iq0";
        pll1_inclk1_logical_to_physical_mapping: string  := "iq1";
        pll1_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll1_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll1_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll1_inclk5_logical_to_physical_mapping: string  := "pld_clk";
        pll1_inclk6_logical_to_physical_mapping: string  := "clkrefclk0";
        pll1_inclk7_logical_to_physical_mapping: string  := "clkrefclk1";
        pll2_inclk0_logical_to_physical_mapping: string  := "iq0";
        pll2_inclk1_logical_to_physical_mapping: string  := "iq1";
        pll2_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll2_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll2_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll2_inclk5_logical_to_physical_mapping: string  := "pld_clk";
        pll2_inclk6_logical_to_physical_mapping: string  := "clkrefclk0";
        pll2_inclk7_logical_to_physical_mapping: string  := "clkrefclk1";
        sim_dump_dprio_internal_reg_at_time: integer := 0;
        sim_dump_filename: string  := "sim_dprio_dump.txt"
    );
    port(
        sync_status     : in     vl_logic_vector(3 downto 0);
        align_status    : in     vl_logic;
        mdio_in         : in     vl_logic;
        mdc             : in     vl_logic;
        port_addr       : in     vl_logic_vector(4 downto 0);
        dev_addr        : in     vl_logic_vector(4 downto 0);
        mdio_dis        : in     vl_logic;
        dprioload       : in     vl_logic;
        mdio_rst        : in     vl_logic;
        cmudividerdprioin: in     vl_logic_vector(29 downto 0);
        cmuplldprioin   : in     vl_logic_vector(119 downto 0);
        cmudprioin      : in     vl_logic_vector(29 downto 0);
        refclkdividerdprioin: in     vl_logic_vector(1 downto 0);
        rxdprioin       : in     vl_logic_vector;
        txdprioin       : in     vl_logic_vector;
        cmudividerdprioout: out    vl_logic_vector(29 downto 0);
        cmuplldprioout  : out    vl_logic_vector(119 downto 0);
        cmudprioout     : out    vl_logic_vector(29 downto 0);
        refclkdividerdprioout: out    vl_logic_vector(1 downto 0);
        rxdprioout      : out    vl_logic_vector;
        txdprioout      : out    vl_logic_vector;
        mdio_out        : out    vl_logic;
        data_enable_n   : out    vl_logic;
        mdio_curr_st    : out    vl_logic_vector(2 downto 0)
    );
end stratixiigx_hssi_cmu_dprio_top;
