library verilog;
use verilog.vl_types.all;
entity \STRATIXII_PRIM_DFFE\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \STRATIXII_PRIM_DFFE\;
