library verilog;
use verilog.vl_types.all;
entity stratixiii_io_ibuf is
    generic(
        differential_mode: string  := "false";
        bus_hold        : string  := "false";
        simulate_z_as   : string  := "Z";
        lpm_type        : string  := "stratixiii_io_ibuf"
    );
    port(
        i               : in     vl_logic;
        ibar            : in     vl_logic;
        dynamicterminationcontrol: in     vl_logic;
        o               : out    vl_logic
    );
end stratixiii_io_ibuf;
