library verilog;
use verilog.vl_types.all;
entity arriaii_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end arriaii_routing_wire;
