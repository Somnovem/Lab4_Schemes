library verilog;
use verilog.vl_types.all;
entity arriaii_hssi_rx_digi_comp_chnl_top is
    port(
        align_status    : in     vl_logic;
        align_status_sync: out    vl_logic;
        align_status_sync_0: in     vl_logic;
        align_status_sync_2: in     vl_logic;
        audi            : in     vl_logic_vector(13 downto 0);
        audi_pre        : in     vl_logic_vector(13 downto 0);
        cg_comp_rd_d_ch0: in     vl_logic;
        cg_comp_rd_d_ch1: in     vl_logic;
        cg_comp_rd_d_ch2: in     vl_logic;
        cg_comp_rd_d_ch3: in     vl_logic;
        cg_comp_rd_d_out: out    vl_logic;
        cg_comp_wr_ch0  : in     vl_logic;
        cg_comp_wr_ch1  : in     vl_logic;
        cg_comp_wr_ch2  : in     vl_logic;
        cg_comp_wr_ch3  : in     vl_logic;
        cg_comp_wr_out  : out    vl_logic;
        clk_1           : in     vl_logic;
        clk_2           : in     vl_logic;
        cmpfifourst     : in     vl_logic;
        comp_curr_st    : out    vl_logic_vector(1 downto 0);
        cudi            : out    vl_logic_vector(31 downto 0);
        cudi_valid      : out    vl_logic;
        del_cond_met_0  : in     vl_logic;
        del_cond_met_out: out    vl_logic;
        dskwclksel      : in     vl_logic_vector(1 downto 0);
        fifo_cnt        : out    vl_logic_vector(4 downto 0);
        fifo_ovr_0      : in     vl_logic;
        fifo_ovr_out    : out    vl_logic;
        fifo_rd_in_comp_0: in     vl_logic;
        fifo_rd_in_comp_2: in     vl_logic;
        fifo_rd_out_comp: out    vl_logic;
        gen2ngen1       : in     vl_logic;
        gen2ngen1_bundle: in     vl_logic;
        hard_reset      : in     vl_logic;
        inferred_rxvalid: in     vl_logic;
        insert_incomplete_0: in     vl_logic;
        insert_incomplete_out: out    vl_logic;
        is_lane0        : in     vl_logic;
        latency_comp_0  : in     vl_logic;
        latency_comp_out: out    vl_logic;
        rauto_speed_ena : in     vl_logic;
        rclkcmpinsertpad: in     vl_logic;
        rclkcmpsq1n     : in     vl_logic_vector(19 downto 0);
        rclkcmpsq1p     : in     vl_logic_vector(19 downto 0);
        rclkcmpsqmd     : in     vl_logic;
        rcmpfifourst    : in     vl_logic;
        rdel_threshold  : in     vl_logic_vector(4 downto 0);
        rdenable        : in     vl_logic;
        rdfifo_almost_empty: out    vl_logic;
        rdfifo_almost_full: out    vl_logic;
        rdfifo_empty    : out    vl_logic;
        rdfifo_full     : out    vl_logic;
        rdwidth_rx      : in     vl_logic;
        rempty_threshold: in     vl_logic_vector(2 downto 0);
        rev_loop_data   : out    vl_logic_vector(19 downto 0);
        rfreq_sel       : in     vl_logic;
        rfull_threshold : in     vl_logic_vector(4 downto 0);
        rgenericfifo    : in     vl_logic;
        rindv_rx        : in     vl_logic;
        rins_threshold  : in     vl_logic_vector(4 downto 0);
        rmatchen        : in     vl_logic;
        rrx_pipe_enable : in     vl_logic;
        rskpsetbased    : in     vl_logic;
        rstart_threshold: in     vl_logic_vector(2 downto 0);
        rtruebac2bac    : in     vl_logic;
        rwa_6g_en       : in     vl_logic;
        scan_mode       : in     vl_logic;
        skpos_det       : out    vl_logic;
        soft_reset      : in     vl_logic;
        sudi            : in     vl_logic_vector(27 downto 0);
        sudi_pre        : in     vl_logic_vector(13 downto 0);
        sync_status     : in     vl_logic;
        wrenable        : in     vl_logic
    );
end arriaii_hssi_rx_digi_comp_chnl_top;
