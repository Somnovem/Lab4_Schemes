library verilog;
use verilog.vl_types.all;
entity cycloneiiils_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end cycloneiiils_routing_wire;
