library verilog;
use verilog.vl_types.all;
entity arriagx_hssi_rx_comp_chnl_top is
    port(
        align_status    : in     vl_logic;
        align_status_sync: out    vl_logic;
        align_status_sync_0: in     vl_logic;
        align_status_sync_2: in     vl_logic;
        audi            : in     vl_logic_vector(13 downto 0);
        audi_pre        : in     vl_logic_vector(13 downto 0);
        clk_1           : in     vl_logic;
        clk_2           : in     vl_logic;
        cmpfifourst     : in     vl_logic;
        comp_curr_st    : out    vl_logic_vector(1 downto 0);
        cudi            : out    vl_logic_vector(31 downto 0);
        cudi_valid      : out    vl_logic;
        disable_fifo_rd : out    vl_logic;
        disable_fifo_rd_0: in     vl_logic;
        disable_fifo_rd_2: in     vl_logic;
        disable_fifo_wr : out    vl_logic;
        disable_fifo_wr_0: in     vl_logic;
        disable_fifo_wr_2: in     vl_logic;
        dskwclksel      : in     vl_logic_vector(1 downto 0);
        fifo_cnt        : out    vl_logic_vector(4 downto 0);
        fifo_rd_in_comp_0: in     vl_logic;
        fifo_rd_in_comp_2: in     vl_logic;
        fifo_rd_out_comp: out    vl_logic;
        hard_reset      : in     vl_logic;
        is_lane0        : in     vl_logic;
        ralempty        : in     vl_logic_vector(3 downto 0);
        ralfull         : in     vl_logic_vector(3 downto 0);
        rclkcmpinsertpad: in     vl_logic;
        rclkcmppos      : in     vl_logic;
        rclkcmpsq1n     : in     vl_logic_vector(19 downto 0);
        rclkcmpsq1p     : in     vl_logic_vector(19 downto 0);
        rclkcmpsqmd     : in     vl_logic;
        rcmpfifourst    : in     vl_logic;
        rdenable        : in     vl_logic;
        rdfifo_almost_empty: out    vl_logic;
        rdfifo_almost_full: out    vl_logic;
        rdfifo_empty    : out    vl_logic;
        rdfifo_full     : out    vl_logic;
        rdwidth_rx      : in     vl_logic;
        rev_loop_data   : out    vl_logic_vector(19 downto 0);
        rgenericfifo    : in     vl_logic;
        rmatchen        : in     vl_logic;
        rrx_pipe_enable : in     vl_logic;
        rskpsetbased    : in     vl_logic;
        rtruebac2bac    : in     vl_logic;
        rwa_6g_en       : in     vl_logic;
        scan_mode       : in     vl_logic;
        soft_reset      : in     vl_logic;
        sudi            : in     vl_logic_vector(27 downto 0);
        sudi_pre        : in     vl_logic_vector(13 downto 0);
        sync_status     : in     vl_logic;
        wrenable        : in     vl_logic
    );
end arriagx_hssi_rx_comp_chnl_top;
