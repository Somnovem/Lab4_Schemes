library verilog;
use verilog.vl_types.all;
entity stratixiigx_hssi_cmu_dprio_reg is
    generic(
        rx_dprio_width  : integer := 800;
        tx_dprio_width  : integer := 400;
        rx0_phy         : integer := 0;
        rx1_phy         : integer := 1;
        rx2_phy         : integer := 2;
        rx3_phy         : integer := 3;
        tx0_phy         : integer := 0;
        tx1_phy         : integer := 1;
        tx2_phy         : integer := 2;
        tx3_phy         : integer := 3;
        rx0_cru_clock0_physical_mapping: string  := "refclk0";
        rx0_cru_clock1_physical_mapping: string  := "refclk1";
        rx0_cru_clock2_physical_mapping: string  := "iq0";
        rx0_cru_clock3_physical_mapping: string  := "iq1";
        rx0_cru_clock4_physical_mapping: string  := "iq2";
        rx0_cru_clock5_physical_mapping: string  := "iq3";
        rx0_cru_clock6_physical_mapping: string  := "iq4";
        rx0_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx0_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        rx1_cru_clock0_physical_mapping: string  := "refclk0";
        rx1_cru_clock1_physical_mapping: string  := "refclk1";
        rx1_cru_clock2_physical_mapping: string  := "iq0";
        rx1_cru_clock3_physical_mapping: string  := "iq1";
        rx1_cru_clock4_physical_mapping: string  := "iq2";
        rx1_cru_clock5_physical_mapping: string  := "iq3";
        rx1_cru_clock6_physical_mapping: string  := "iq4";
        rx1_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx1_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        rx2_cru_clock0_physical_mapping: string  := "refclk0";
        rx2_cru_clock1_physical_mapping: string  := "refclk1";
        rx2_cru_clock2_physical_mapping: string  := "iq0";
        rx2_cru_clock3_physical_mapping: string  := "iq1";
        rx2_cru_clock4_physical_mapping: string  := "iq2";
        rx2_cru_clock5_physical_mapping: string  := "iq3";
        rx2_cru_clock6_physical_mapping: string  := "iq4";
        rx2_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx2_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        rx3_cru_clock0_physical_mapping: string  := "refclk0";
        rx3_cru_clock1_physical_mapping: string  := "refclk1";
        rx3_cru_clock2_physical_mapping: string  := "iq0";
        rx3_cru_clock3_physical_mapping: string  := "iq1";
        rx3_cru_clock4_physical_mapping: string  := "iq2";
        rx3_cru_clock5_physical_mapping: string  := "iq3";
        rx3_cru_clock6_physical_mapping: string  := "iq4";
        rx3_cru_clock7_physical_mapping: string  := "pld_cru_clk";
        rx3_cru_clock8_physical_mapping: string  := "cmu_div_clk";
        tx0_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx0_pll_fast_clk1_physical_mapping: string  := "pll1";
        tx1_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx1_pll_fast_clk1_physical_mapping: string  := "pll1";
        tx2_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx2_pll_fast_clk1_physical_mapping: string  := "pll1";
        tx3_pll_fast_clk0_physical_mapping: string  := "pll0";
        tx3_pll_fast_clk1_physical_mapping: string  := "pll1";
        pll0_phy        : integer := 0;
        pll1_phy        : integer := 1;
        pll2_phy        : integer := 2;
        pll0_inclk0_logical_to_physical_mapping: string  := "iq0";
        pll0_inclk1_logical_to_physical_mapping: string  := "iq1";
        pll0_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll0_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll0_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll0_inclk5_logical_to_physical_mapping: string  := "pld_clk";
        pll0_inclk6_logical_to_physical_mapping: string  := "clkrefclk0";
        pll0_inclk7_logical_to_physical_mapping: string  := "clkrefclk1";
        pll1_inclk0_logical_to_physical_mapping: string  := "iq0";
        pll1_inclk1_logical_to_physical_mapping: string  := "iq1";
        pll1_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll1_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll1_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll1_inclk5_logical_to_physical_mapping: string  := "pld_clk";
        pll1_inclk6_logical_to_physical_mapping: string  := "clkrefclk0";
        pll1_inclk7_logical_to_physical_mapping: string  := "clkrefclk1";
        pll2_inclk0_logical_to_physical_mapping: string  := "iq0";
        pll2_inclk1_logical_to_physical_mapping: string  := "iq1";
        pll2_inclk2_logical_to_physical_mapping: string  := "iq2";
        pll2_inclk3_logical_to_physical_mapping: string  := "iq3";
        pll2_inclk4_logical_to_physical_mapping: string  := "iq4";
        pll2_inclk5_logical_to_physical_mapping: string  := "pld_clk";
        pll2_inclk6_logical_to_physical_mapping: string  := "clkrefclk0";
        pll2_inclk7_logical_to_physical_mapping: string  := "clkrefclk1";
        sim_dump_dprio_internal_reg_at_time: integer := 0;
        sim_dump_filename: string  := "sim_dprio_dump.txt";
        \XGXS_CTRL\     : integer := 0;
        \XGXS_STATUS1\  : integer := 1;
        \XGXS_STATUS2\  : integer := 8;
        \XGXS_LANE_STATUS\: integer := 24;
        \TRUNKING_MODE\ : integer := 32768;
        \PCS_CTRL1_CH0\ : integer := 32769;
        \PCS_CTRL1_CH1\ : integer := 32770;
        \PCS_CTRL1_CH2\ : integer := 32771;
        \PCS_CTRL1_CH3\ : integer := 32772;
        \PCS_CTRL2_CH0\ : integer := 32773;
        \PCS_CTRL2_CH1\ : integer := 32774;
        \PCS_CTRL2_CH2\ : integer := 32775;
        \PCS_CTRL2_CH3\ : integer := 32776;
        \PCS_CTRL3_CH0\ : integer := 32777;
        \PCS_CTRL3_CH1\ : integer := 32778;
        \PCS_CTRL3_CH2\ : integer := 32779;
        \PCS_CTRL3_CH3\ : integer := 32780;
        \PCS_CTRL4_CH0\ : integer := 32781;
        \PCS_CTRL4_CH1\ : integer := 32782;
        \PCS_CTRL4_CH2\ : integer := 32783;
        \PCS_CTRL4_CH3\ : integer := 32784;
        \PCS_CTRL5_CH0\ : integer := 32785;
        \PCS_CTRL5_CH1\ : integer := 32786;
        \PCS_CTRL5_CH2\ : integer := 32787;
        \PCS_CTRL5_CH3\ : integer := 32788;
        \PCS_CTRL6_CH0\ : integer := 32789;
        \PCS_CTRL6_CH1\ : integer := 32790;
        \PCS_CTRL6_CH2\ : integer := 32791;
        \PCS_CTRL6_CH3\ : integer := 32792;
        \PCS_CTRL7_CH0\ : integer := 32793;
        \PCS_CTRL7_CH1\ : integer := 32794;
        \PCS_CTRL7_CH2\ : integer := 32795;
        \PCS_CTRL7_CH3\ : integer := 32796;
        \PCS_CTRL8_CH0\ : integer := 32797;
        \PCS_CTRL8_CH1\ : integer := 32798;
        \PCS_CTRL8_CH2\ : integer := 32799;
        \PCS_CTRL8_CH3\ : integer := 32800;
        \PRBS_BIST_CTRL_CH0\: integer := 32801;
        \PRBS_BIST_CTRL_CH1\: integer := 32802;
        \PRBS_BIST_CTRL_CH2\: integer := 32803;
        \PRBS_BIST_CTRL_CH3\: integer := 32804;
        \PCS_CTRL9_CH0\ : integer := 32805;
        \PCS_CTRL9_CH1\ : integer := 32806;
        \PCS_CTRL9_CH2\ : integer := 32807;
        \PCS_CTRL9_CH3\ : integer := 32808;
        \PCS_CTRL10_CH0\: integer := 32809;
        \PCS_CTRL10_CH1\: integer := 32810;
        \PCS_CTRL10_CH2\: integer := 32811;
        \PCS_CTRL10_CH3\: integer := 32812;
        \PCS_CTRL11_CH0\: integer := 32813;
        \PCS_CTRL11_CH1\: integer := 32814;
        \PCS_CTRL11_CH2\: integer := 32815;
        \PCS_CTRL11_CH3\: integer := 32816;
        \PCS_CTRL12_CH0\: integer := 32817;
        \PCS_CTRL12_CH1\: integer := 32818;
        \PCS_CTRL12_CH2\: integer := 32819;
        \PCS_CTRL12_CH3\: integer := 32820;
        \PCS_CTRL13_CH0\: integer := 32821;
        \PCS_CTRL13_CH1\: integer := 32822;
        \PCS_CTRL13_CH2\: integer := 32823;
        \PCS_CTRL13_CH3\: integer := 32824;
        \PCS_CTRL14_CH0\: integer := 32825;
        \PCS_CTRL14_CH1\: integer := 32826;
        \PCS_CTRL14_CH2\: integer := 32827;
        \PCS_CTRL14_CH3\: integer := 32828;
        \PCS_CTRL15_CH0\: integer := 32829;
        \PCS_CTRL15_CH1\: integer := 32830;
        \PCS_CTRL15_CH2\: integer := 32831;
        \PCS_CTRL15_CH3\: integer := 32832;
        \PCS_GLOBAL_CTRL0\: integer := 32848;
        \PCS_GLOBAL_CTRL1\: integer := 32849;
        \PCS_GLOBAL_CTRL2\: integer := 32850;
        \PMA_CTRL1_CH0\ : integer := 32864;
        \PMA_CTRL1_CH1\ : integer := 32865;
        \PMA_CTRL1_CH2\ : integer := 32866;
        \PMA_CTRL1_CH3\ : integer := 32867;
        \PMA_CTRL2_CH0\ : integer := 32868;
        \PMA_CTRL2_CH1\ : integer := 32869;
        \PMA_CTRL2_CH2\ : integer := 32870;
        \PMA_CTRL2_CH3\ : integer := 32871;
        \PMA_CTRL3_CH0\ : integer := 32872;
        \PMA_CTRL3_CH1\ : integer := 32873;
        \PMA_CTRL3_CH2\ : integer := 32874;
        \PMA_CTRL3_CH3\ : integer := 32875;
        \PMA_CTRL4_CH0\ : integer := 32876;
        \PMA_CTRL4_CH1\ : integer := 32877;
        \PMA_CTRL4_CH2\ : integer := 32878;
        \PMA_CTRL4_CH3\ : integer := 32879;
        \PMA_CTRL5_CH0\ : integer := 32880;
        \PMA_CTRL5_CH1\ : integer := 32881;
        \PMA_CTRL5_CH2\ : integer := 32882;
        \PMA_CTRL5_CH3\ : integer := 32883;
        \PMA_CTRL6_CH0\ : integer := 32884;
        \PMA_CTRL6_CH1\ : integer := 32885;
        \PMA_CTRL6_CH2\ : integer := 32886;
        \PMA_CTRL6_CH3\ : integer := 32887;
        \PMA_CTRL7_CH0\ : integer := 32888;
        \PMA_CTRL7_CH1\ : integer := 32889;
        \PMA_CTRL7_CH2\ : integer := 32890;
        \PMA_CTRL7_CH3\ : integer := 32891;
        \PMA_CTRL8_CH0\ : integer := 32892;
        \PMA_CTRL8_CH1\ : integer := 32893;
        \PMA_CTRL8_CH2\ : integer := 32894;
        \PMA_CTRL8_CH3\ : integer := 32895;
        \PMA_CTRL9_CH0\ : integer := 32896;
        \PMA_CTRL9_CH1\ : integer := 32897;
        \PMA_CTRL9_CH2\ : integer := 32898;
        \PMA_CTRL9_CH3\ : integer := 32899;
        \PMA_CTRL10_CH0\: integer := 32900;
        \PMA_CTRL10_CH1\: integer := 32901;
        \PMA_CTRL10_CH2\: integer := 32902;
        \PMA_CTRL10_CH3\: integer := 32903;
        \PMA_CTRL11_CH0\: integer := 32904;
        \PMA_CTRL11_CH1\: integer := 32905;
        \PMA_CTRL11_CH2\: integer := 32906;
        \PMA_CTRL11_CH3\: integer := 32907;
        \PMA_GLOBAL_CTRL0\: integer := 32912;
        \PMA_GLOBAL_CTRL1\: integer := 32913;
        \PMA_GLOBAL_CTRL2\: integer := 32914;
        \PMA_GLOBAL_CTRL3\: integer := 32915;
        \PMA_GLOBAL_CTRL4\: integer := 32916;
        \PMA_GLOBAL_CTRL5\: integer := 32917;
        \PMA_GLOBAL_CTRL6\: integer := 32918;
        \PMA_GLOBAL_CTRL7\: integer := 32919;
        \PMA_GLOBAL_CTRL8\: integer := 32920;
        \PMA_GLOBAL_CTRL9\: integer := 32921
    );
    port(
        mdc             : in     vl_logic;
        mdio_rst        : in     vl_logic;
        mdio_dis        : in     vl_logic;
        dprioload       : in     vl_logic;
        align_status    : in     vl_logic;
        sync_status     : in     vl_logic_vector(3 downto 0);
        reg_addr        : in     vl_logic_vector(15 downto 0);
        mdio_wr         : in     vl_logic;
        mdio_rd         : in     vl_logic;
        dev_addr_0      : in     vl_logic;
        mbus_in         : in     vl_logic_vector(15 downto 0);
        cmudividerdprioin: in     vl_logic_vector(29 downto 0);
        cmuplldprioin   : in     vl_logic_vector(119 downto 0);
        cmudprioin      : in     vl_logic_vector(29 downto 0);
        refclkdividerdprioin: in     vl_logic_vector(1 downto 0);
        rxdprioin       : in     vl_logic_vector;
        txdprioin       : in     vl_logic_vector;
        cmudividerdprioout: out    vl_logic_vector(29 downto 0);
        cmuplldprioout  : out    vl_logic_vector(119 downto 0);
        cmudprioout     : out    vl_logic_vector(29 downto 0);
        refclkdividerdprioout: out    vl_logic_vector(1 downto 0);
        rxdprioout      : out    vl_logic_vector;
        txdprioout      : out    vl_logic_vector;
        mbus_out        : out    vl_logic_vector(15 downto 0)
    );
end stratixiigx_hssi_cmu_dprio_reg;
