library verilog;
use verilog.vl_types.all;
entity arriagx_hssi_tx_digi is
    port(
        txpcs_rst       : in     vl_logic;
        scan_mode       : in     vl_logic;
        txd             : in     vl_logic_vector(43 downto 0);
        pld_tx_clk      : in     vl_logic;
        polinv_tx       : in     vl_logic;
        rev_loop_data   : in     vl_logic_vector(19 downto 0);
        wrenable_tx     : in     vl_logic;
        rddisable_tx    : in     vl_logic;
        phfifourst_tx   : in     vl_logic;
        txfifo_shared_sig_in_ch0: in     vl_logic_vector(3 downto 0);
        txfifo_shared_sig_in_q0_ch0: in     vl_logic_vector(3 downto 0);
        txfifo_shared_sig_out: out    vl_logic_vector(3 downto 0);
        full_tx         : out    vl_logic;
        empty_tx        : out    vl_logic;
        tx_data_ts      : in     vl_logic_vector(7 downto 0);
        tx_ctl_ts       : in     vl_logic;
        refclk_pma      : in     vl_logic;
        txpma_local_clk : in     vl_logic;
        tx_clk_out      : out    vl_logic;
        tx_data_tc      : out    vl_logic_vector(7 downto 0);
        tx_ctl_tc       : out    vl_logic;
        pudr            : out    vl_logic_vector(19 downto 0);
        rd_enable_sync  : out    vl_logic;
        refclk_b        : out    vl_logic;
        txlp20b         : out    vl_logic_vector(19 downto 0);
        tx_pipe_clk     : out    vl_logic;
        encoder_testbus : out    vl_logic_vector(9 downto 0);
        tx_ctrl_testbus : out    vl_logic_vector(9 downto 0);
        tx_pipe_soft_reset: out    vl_logic;
        tx_pipe_electidle: out    vl_logic;
        rrev_loopbk     : in     vl_logic;
        rev_loopbk      : in     vl_logic;
        rbisten_tx      : in     vl_logic;
        rforce_disp     : in     vl_logic;
        rib_force_disp  : in     vl_logic;
        rforce_echar    : in     vl_logic;
        rforce_kchar    : in     vl_logic;
        rendec_tx       : in     vl_logic;
        rge_xaui_tx     : in     vl_logic;
        rdwidth_tx      : in     vl_logic;
        rtxfifo_dis     : in     vl_logic;
        rcascaded_8b10b_en_tx: in     vl_logic;
        rprbsen_tx      : in     vl_logic;
        rprbs_sel       : in     vl_logic_vector(2 downto 0);
        rbist_sel       : in     vl_logic_vector(1 downto 0);
        rcxpat_chnl_en  : in     vl_logic_vector(1 downto 0);
        renpolinv_tx    : in     vl_logic;
        rphfifopldentx  : in     vl_logic;
        rphfifoursttx   : in     vl_logic;
        rfreerun_tx     : in     vl_logic;
        rtxwrclksel     : in     vl_logic;
        rtxrdclksel     : in     vl_logic;
        renbitrev_tx    : in     vl_logic;
        rensymswap_tx   : in     vl_logic;
        r8b10b_enc_ibm_en: in     vl_logic;
        rtxfifo_lowlatency_en: in     vl_logic;
        rpmadwidth_tx   : in     vl_logic;
        rpma_doublewidth_tx: in     vl_logic;
        rtx_pipe_enable : in     vl_logic;
        rindv_tx        : in     vl_logic;
        rendec_data_sel_tx: in     vl_logic;
        rphfifo_master_sel_tx: in     vl_logic
    );
end arriagx_hssi_tx_digi;
