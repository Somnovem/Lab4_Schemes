library verilog;
use verilog.vl_types.all;
entity stratixiv_hssi_pma_c_rx is
    generic(
        \PARAM_DELAY\   : integer := 0;
        \SD_PULSE_DELAY\: integer := 1;
        \INVALID_SD_ON_OFF\: integer := 500
    );
    port(
        ac_mode         : in     vl_logic;
        analog_sd       : out    vl_logic;
        atb0_rx         : inout  vl_logic;
        atb1_rx         : inout  vl_logic;
        atbsel          : in     vl_logic_vector(5 downto 0);
        bsmode          : in     vl_logic;
        bsrxn_in        : in     vl_logic;
        bsrxn_out       : out    vl_logic;
        bsrxp_in        : in     vl_logic;
        bsrxp_out       : out    vl_logic;
        ck0_sigdet      : in     vl_logic;
        eqa_ctrl        : in     vl_logic;
        eqb_ctrl        : in     vl_logic;
        eqc_ctrl        : in     vl_logic;
        eqd_ctrl        : in     vl_logic;
        eqv_ctrl        : inout  vl_logic;
        ibc50u          : inout  vl_logic_vector(1 downto 0);
        ibp50u          : inout  vl_logic_vector(3 downto 0);
        ibp150u         : inout  vl_logic_vector(1 downto 0);
        inn             : inout  vl_logic;
        inn3            : out    vl_logic;
        inp             : inout  vl_logic;
        inp3            : out    vl_logic;
        lpbkn           : in     vl_logic;
        lpbkp           : in     vl_logic;
        mem_init        : in     vl_logic;
        oc_calpd        : in     vl_logic;
        oc_en           : in     vl_logic;
        pd2             : out    vl_logic;
        pd2_term        : in     vl_logic;
        pd_rxclk_term   : out    vl_logic;
        pdb             : in     vl_logic;
        pdb_clk         : in     vl_logic;
        pdbh_rx         : out    vl_logic;
        pdbh_rxclk_term : out    vl_logic;
        pdbh_term       : in     vl_logic;
        pdshft_clk      : in     vl_logic;
        rbit_dc         : in     vl_logic_vector(3 downto 0);
        rdlpbkn         : out    vl_logic;
        rdlpbkn_far     : out    vl_logic;
        rdlpbkp         : out    vl_logic;
        rdlpbkp_far     : out    vl_logic;
        refclk          : in     vl_logic;
        rstn            : in     vl_logic;
        rx_b50          : in     vl_logic_vector(3 downto 0);
        rx_oc           : in     vl_logic_vector(7 downto 0);
        rx_test         : in     vl_logic;
        rx_testclk      : in     vl_logic;
        rxbuf_ibias     : out    vl_logic;
        rxn             : out    vl_logic;
        rxp             : out    vl_logic;
        s_lpbk          : in     vl_logic;
        s_rdlpbk        : in     vl_logic;
        sd_cdr          : out    vl_logic;
        sd_cpon         : out    vl_logic;
        sd_cpop         : out    vl_logic;
        sd_force        : in     vl_logic;
        sd_off          : in     vl_logic_vector(4 downto 0);
        sd_on           : in     vl_logic_vector(3 downto 0);
        sdlv            : in     vl_logic_vector(3 downto 0);
        slew            : in     vl_logic_vector(1 downto 0);
        term            : in     vl_logic_vector(2 downto 0);
        vcce_la         : in     vl_logic;
        vcce_oa         : in     vl_logic;
        vccehtxqyx      : in     vl_logic;
        vssexqyx        : in     vl_logic;
        vtt             : in     vl_logic_vector(2 downto 0)
    );
end stratixiv_hssi_pma_c_rx;
