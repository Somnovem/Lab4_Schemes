library verilog;
use verilog.vl_types.all;
entity \ALTERA_MF_MEMORY_INITIALIZATION\ is
end \ALTERA_MF_MEMORY_INITIALIZATION\;
