library verilog;
use verilog.vl_types.all;
entity \STRATIX_PRIM_DFFEAS\ is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end \STRATIX_PRIM_DFFEAS\;
